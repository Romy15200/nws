/*
*
*	Taken from VIS Benchmarks <ftp://vlsi.colorado.edu/pub/vis/vis-verilog-models-1.3.tar.gz>
*	Modified by Ahmed Irfan <irfan@fbk.eu>
*
*/
//Author: Fabio Somenzi <Fabio@Colorado.EDU>
// Slider puzzle with N rows and N columns.             +-------+----+----+----+-----+-----+
//                                                      |  0    |  1 |  2 |  3 |.....| N-1 |
// The entries of the matrix are numbered thus:         +-------+----+----+----+-----+-----+
//                                                      |  N    | N+1| N+2| N+3|.....| 2N-1|
//                                                      +-------+----+----+----+-----+-----+  
//                                                      |.......|....|....|....|.....|.....|          
//                                                      +-------+----+----+----+-----+-----+
//                                                      |(N-1)*N|....|....|....|.....|N^2-1|
//                                                      +-------+----+----+----+-----+-----+
module slidingBoard(clock,from,to);
    input       clock;
    input [15:0] from;
    input [15:0] to;

    reg [15:0] 	b[0:65535];
    reg [15:0] 	freg, treg;
    wire 	valid, parity;

    initial begin
        for (i=0; i < 65536; i = i+1) begin
          b[i] = 65535-i;
	end
        treg = 0;
	freg = 0;
    end 

    assign valid = (b[treg] == 16'b0) &&
                    ( //sliding between rows
		   (treg[5:0] == freg[5:0] && ((freg[15:8] == 0 && treg[15:8] == 1) || 
(treg[15:8] == 0 && freg[15:8] == 1) || 
(freg[15:8] == 1 && treg[15:8] == 2) || 
(treg[15:8] == 1 && freg[15:8] == 2) || 
(freg[15:8] == 2 && treg[15:8] == 3) || 
(treg[15:8] == 2 && freg[15:8] == 3) || 
(freg[15:8] == 3 && treg[15:8] == 4) || 
(treg[15:8] == 3 && freg[15:8] == 4) || 
(freg[15:8] == 4 && treg[15:8] == 5) || 
(treg[15:8] == 4 && freg[15:8] == 5) || 
(freg[15:8] == 5 && treg[15:8] == 6) || 
(treg[15:8] == 5 && freg[15:8] == 6) || 
(freg[15:8] == 6 && treg[15:8] == 7) || 
(treg[15:8] == 6 && freg[15:8] == 7) || 
(freg[15:8] == 7 && treg[15:8] == 8) || 
(treg[15:8] == 7 && freg[15:8] == 8) || 
(freg[15:8] == 8 && treg[15:8] == 9) || 
(treg[15:8] == 8 && freg[15:8] == 9) || 
(freg[15:8] == 9 && treg[15:8] == 10) || 
(treg[15:8] == 9 && freg[15:8] == 10) || 
(freg[15:8] == 10 && treg[15:8] == 11) || 
(treg[15:8] == 10 && freg[15:8] == 11) || 
(freg[15:8] == 11 && treg[15:8] == 12) || 
(treg[15:8] == 11 && freg[15:8] == 12) || 
(freg[15:8] == 12 && treg[15:8] == 13) || 
(treg[15:8] == 12 && freg[15:8] == 13) || 
(freg[15:8] == 13 && treg[15:8] == 14) || 
(treg[15:8] == 13 && freg[15:8] == 14) || 
(freg[15:8] == 14 && treg[15:8] == 15) || 
(treg[15:8] == 14 && freg[15:8] == 15) || 
(freg[15:8] == 15 && treg[15:8] == 16) || 
(treg[15:8] == 15 && freg[15:8] == 16) || 
(freg[15:8] == 16 && treg[15:8] == 17) || 
(treg[15:8] == 16 && freg[15:8] == 17) || 
(freg[15:8] == 17 && treg[15:8] == 18) || 
(treg[15:8] == 17 && freg[15:8] == 18) || 
(freg[15:8] == 18 && treg[15:8] == 19) || 
(treg[15:8] == 18 && freg[15:8] == 19) || 
(freg[15:8] == 19 && treg[15:8] == 20) || 
(treg[15:8] == 19 && freg[15:8] == 20) || 
(freg[15:8] == 20 && treg[15:8] == 21) || 
(treg[15:8] == 20 && freg[15:8] == 21) || 
(freg[15:8] == 21 && treg[15:8] == 22) || 
(treg[15:8] == 21 && freg[15:8] == 22) || 
(freg[15:8] == 22 && treg[15:8] == 23) || 
(treg[15:8] == 22 && freg[15:8] == 23) || 
(freg[15:8] == 23 && treg[15:8] == 24) || 
(treg[15:8] == 23 && freg[15:8] == 24) || 
(freg[15:8] == 24 && treg[15:8] == 25) || 
(treg[15:8] == 24 && freg[15:8] == 25) || 
(freg[15:8] == 25 && treg[15:8] == 26) || 
(treg[15:8] == 25 && freg[15:8] == 26) || 
(freg[15:8] == 26 && treg[15:8] == 27) || 
(treg[15:8] == 26 && freg[15:8] == 27) || 
(freg[15:8] == 27 && treg[15:8] == 28) || 
(treg[15:8] == 27 && freg[15:8] == 28) || 
(freg[15:8] == 28 && treg[15:8] == 29) || 
(treg[15:8] == 28 && freg[15:8] == 29) || 
(freg[15:8] == 29 && treg[15:8] == 30) || 
(treg[15:8] == 29 && freg[15:8] == 30) || 
(freg[15:8] == 30 && treg[15:8] == 31) || 
(treg[15:8] == 30 && freg[15:8] == 31) || 
(freg[15:8] == 31 && treg[15:8] == 32) || 
(treg[15:8] == 31 && freg[15:8] == 32) || 
(freg[15:8] == 32 && treg[15:8] == 33) || 
(treg[15:8] == 32 && freg[15:8] == 33) || 
(freg[15:8] == 33 && treg[15:8] == 34) || 
(treg[15:8] == 33 && freg[15:8] == 34) || 
(freg[15:8] == 34 && treg[15:8] == 35) || 
(treg[15:8] == 34 && freg[15:8] == 35) || 
(freg[15:8] == 35 && treg[15:8] == 36) || 
(treg[15:8] == 35 && freg[15:8] == 36) || 
(freg[15:8] == 36 && treg[15:8] == 37) || 
(treg[15:8] == 36 && freg[15:8] == 37) || 
(freg[15:8] == 37 && treg[15:8] == 38) || 
(treg[15:8] == 37 && freg[15:8] == 38) || 
(freg[15:8] == 38 && treg[15:8] == 39) || 
(treg[15:8] == 38 && freg[15:8] == 39) || 
(freg[15:8] == 39 && treg[15:8] == 40) || 
(treg[15:8] == 39 && freg[15:8] == 40) || 
(freg[15:8] == 40 && treg[15:8] == 41) || 
(treg[15:8] == 40 && freg[15:8] == 41) || 
(freg[15:8] == 41 && treg[15:8] == 42) || 
(treg[15:8] == 41 && freg[15:8] == 42) || 
(freg[15:8] == 42 && treg[15:8] == 43) || 
(treg[15:8] == 42 && freg[15:8] == 43) || 
(freg[15:8] == 43 && treg[15:8] == 44) || 
(treg[15:8] == 43 && freg[15:8] == 44) || 
(freg[15:8] == 44 && treg[15:8] == 45) || 
(treg[15:8] == 44 && freg[15:8] == 45) || 
(freg[15:8] == 45 && treg[15:8] == 46) || 
(treg[15:8] == 45 && freg[15:8] == 46) || 
(freg[15:8] == 46 && treg[15:8] == 47) || 
(treg[15:8] == 46 && freg[15:8] == 47) || 
(freg[15:8] == 47 && treg[15:8] == 48) || 
(treg[15:8] == 47 && freg[15:8] == 48) || 
(freg[15:8] == 48 && treg[15:8] == 49) || 
(treg[15:8] == 48 && freg[15:8] == 49) || 
(freg[15:8] == 49 && treg[15:8] == 50) || 
(treg[15:8] == 49 && freg[15:8] == 50) || 
(freg[15:8] == 50 && treg[15:8] == 51) || 
(treg[15:8] == 50 && freg[15:8] == 51) || 
(freg[15:8] == 51 && treg[15:8] == 52) || 
(treg[15:8] == 51 && freg[15:8] == 52) || 
(freg[15:8] == 52 && treg[15:8] == 53) || 
(treg[15:8] == 52 && freg[15:8] == 53) || 
(freg[15:8] == 53 && treg[15:8] == 54) || 
(treg[15:8] == 53 && freg[15:8] == 54) || 
(freg[15:8] == 54 && treg[15:8] == 55) || 
(treg[15:8] == 54 && freg[15:8] == 55) || 
(freg[15:8] == 55 && treg[15:8] == 56) || 
(treg[15:8] == 55 && freg[15:8] == 56) || 
(freg[15:8] == 56 && treg[15:8] == 57) || 
(treg[15:8] == 56 && freg[15:8] == 57) || 
(freg[15:8] == 57 && treg[15:8] == 58) || 
(treg[15:8] == 57 && freg[15:8] == 58) || 
(freg[15:8] == 58 && treg[15:8] == 59) || 
(treg[15:8] == 58 && freg[15:8] == 59) || 
(freg[15:8] == 59 && treg[15:8] == 60) || 
(treg[15:8] == 59 && freg[15:8] == 60) || 
(freg[15:8] == 60 && treg[15:8] == 61) || 
(treg[15:8] == 60 && freg[15:8] == 61) || 
(freg[15:8] == 61 && treg[15:8] == 62) || 
(treg[15:8] == 61 && freg[15:8] == 62) || 
(freg[15:8] == 62 && treg[15:8] == 63) || 
(treg[15:8] == 62 && freg[15:8] == 63) || 
(freg[15:8] == 63 && treg[15:8] == 64) || 
(treg[15:8] == 63 && freg[15:8] == 64) || 
(freg[15:8] == 64 && treg[15:8] == 65) || 
(treg[15:8] == 64 && freg[15:8] == 65) || 
(freg[15:8] == 65 && treg[15:8] == 66) || 
(treg[15:8] == 65 && freg[15:8] == 66) || 
(freg[15:8] == 66 && treg[15:8] == 67) || 
(treg[15:8] == 66 && freg[15:8] == 67) || 
(freg[15:8] == 67 && treg[15:8] == 68) || 
(treg[15:8] == 67 && freg[15:8] == 68) || 
(freg[15:8] == 68 && treg[15:8] == 69) || 
(treg[15:8] == 68 && freg[15:8] == 69) || 
(freg[15:8] == 69 && treg[15:8] == 70) || 
(treg[15:8] == 69 && freg[15:8] == 70) || 
(freg[15:8] == 70 && treg[15:8] == 71) || 
(treg[15:8] == 70 && freg[15:8] == 71) || 
(freg[15:8] == 71 && treg[15:8] == 72) || 
(treg[15:8] == 71 && freg[15:8] == 72) || 
(freg[15:8] == 72 && treg[15:8] == 73) || 
(treg[15:8] == 72 && freg[15:8] == 73) || 
(freg[15:8] == 73 && treg[15:8] == 74) || 
(treg[15:8] == 73 && freg[15:8] == 74) || 
(freg[15:8] == 74 && treg[15:8] == 75) || 
(treg[15:8] == 74 && freg[15:8] == 75) || 
(freg[15:8] == 75 && treg[15:8] == 76) || 
(treg[15:8] == 75 && freg[15:8] == 76) || 
(freg[15:8] == 76 && treg[15:8] == 77) || 
(treg[15:8] == 76 && freg[15:8] == 77) || 
(freg[15:8] == 77 && treg[15:8] == 78) || 
(treg[15:8] == 77 && freg[15:8] == 78) || 
(freg[15:8] == 78 && treg[15:8] == 79) || 
(treg[15:8] == 78 && freg[15:8] == 79) || 
(freg[15:8] == 79 && treg[15:8] == 80) || 
(treg[15:8] == 79 && freg[15:8] == 80) || 
(freg[15:8] == 80 && treg[15:8] == 81) || 
(treg[15:8] == 80 && freg[15:8] == 81) || 
(freg[15:8] == 81 && treg[15:8] == 82) || 
(treg[15:8] == 81 && freg[15:8] == 82) || 
(freg[15:8] == 82 && treg[15:8] == 83) || 
(treg[15:8] == 82 && freg[15:8] == 83) || 
(freg[15:8] == 83 && treg[15:8] == 84) || 
(treg[15:8] == 83 && freg[15:8] == 84) || 
(freg[15:8] == 84 && treg[15:8] == 85) || 
(treg[15:8] == 84 && freg[15:8] == 85) || 
(freg[15:8] == 85 && treg[15:8] == 86) || 
(treg[15:8] == 85 && freg[15:8] == 86) || 
(freg[15:8] == 86 && treg[15:8] == 87) || 
(treg[15:8] == 86 && freg[15:8] == 87) || 
(freg[15:8] == 87 && treg[15:8] == 88) || 
(treg[15:8] == 87 && freg[15:8] == 88) || 
(freg[15:8] == 88 && treg[15:8] == 89) || 
(treg[15:8] == 88 && freg[15:8] == 89) || 
(freg[15:8] == 89 && treg[15:8] == 90) || 
(treg[15:8] == 89 && freg[15:8] == 90) || 
(freg[15:8] == 90 && treg[15:8] == 91) || 
(treg[15:8] == 90 && freg[15:8] == 91) || 
(freg[15:8] == 91 && treg[15:8] == 92) || 
(treg[15:8] == 91 && freg[15:8] == 92) || 
(freg[15:8] == 92 && treg[15:8] == 93) || 
(treg[15:8] == 92 && freg[15:8] == 93) || 
(freg[15:8] == 93 && treg[15:8] == 94) || 
(treg[15:8] == 93 && freg[15:8] == 94) || 
(freg[15:8] == 94 && treg[15:8] == 95) || 
(treg[15:8] == 94 && freg[15:8] == 95) || 
(freg[15:8] == 95 && treg[15:8] == 96) || 
(treg[15:8] == 95 && freg[15:8] == 96) || 
(freg[15:8] == 96 && treg[15:8] == 97) || 
(treg[15:8] == 96 && freg[15:8] == 97) || 
(freg[15:8] == 97 && treg[15:8] == 98) || 
(treg[15:8] == 97 && freg[15:8] == 98) || 
(freg[15:8] == 98 && treg[15:8] == 99) || 
(treg[15:8] == 98 && freg[15:8] == 99) || 
(freg[15:8] == 99 && treg[15:8] == 100) || 
(treg[15:8] == 99 && freg[15:8] == 100) || 
(freg[15:8] == 100 && treg[15:8] == 101) || 
(treg[15:8] == 100 && freg[15:8] == 101) || 
(freg[15:8] == 101 && treg[15:8] == 102) || 
(treg[15:8] == 101 && freg[15:8] == 102) || 
(freg[15:8] == 102 && treg[15:8] == 103) || 
(treg[15:8] == 102 && freg[15:8] == 103) || 
(freg[15:8] == 103 && treg[15:8] == 104) || 
(treg[15:8] == 103 && freg[15:8] == 104) || 
(freg[15:8] == 104 && treg[15:8] == 105) || 
(treg[15:8] == 104 && freg[15:8] == 105) || 
(freg[15:8] == 105 && treg[15:8] == 106) || 
(treg[15:8] == 105 && freg[15:8] == 106) || 
(freg[15:8] == 106 && treg[15:8] == 107) || 
(treg[15:8] == 106 && freg[15:8] == 107) || 
(freg[15:8] == 107 && treg[15:8] == 108) || 
(treg[15:8] == 107 && freg[15:8] == 108) || 
(freg[15:8] == 108 && treg[15:8] == 109) || 
(treg[15:8] == 108 && freg[15:8] == 109) || 
(freg[15:8] == 109 && treg[15:8] == 110) || 
(treg[15:8] == 109 && freg[15:8] == 110) || 
(freg[15:8] == 110 && treg[15:8] == 111) || 
(treg[15:8] == 110 && freg[15:8] == 111) || 
(freg[15:8] == 111 && treg[15:8] == 112) || 
(treg[15:8] == 111 && freg[15:8] == 112) || 
(freg[15:8] == 112 && treg[15:8] == 113) || 
(treg[15:8] == 112 && freg[15:8] == 113) || 
(freg[15:8] == 113 && treg[15:8] == 114) || 
(treg[15:8] == 113 && freg[15:8] == 114) || 
(freg[15:8] == 114 && treg[15:8] == 115) || 
(treg[15:8] == 114 && freg[15:8] == 115) || 
(freg[15:8] == 115 && treg[15:8] == 116) || 
(treg[15:8] == 115 && freg[15:8] == 116) || 
(freg[15:8] == 116 && treg[15:8] == 117) || 
(treg[15:8] == 116 && freg[15:8] == 117) || 
(freg[15:8] == 117 && treg[15:8] == 118) || 
(treg[15:8] == 117 && freg[15:8] == 118) || 
(freg[15:8] == 118 && treg[15:8] == 119) || 
(treg[15:8] == 118 && freg[15:8] == 119) || 
(freg[15:8] == 119 && treg[15:8] == 120) || 
(treg[15:8] == 119 && freg[15:8] == 120) || 
(freg[15:8] == 120 && treg[15:8] == 121) || 
(treg[15:8] == 120 && freg[15:8] == 121) || 
(freg[15:8] == 121 && treg[15:8] == 122) || 
(treg[15:8] == 121 && freg[15:8] == 122) || 
(freg[15:8] == 122 && treg[15:8] == 123) || 
(treg[15:8] == 122 && freg[15:8] == 123) || 
(freg[15:8] == 123 && treg[15:8] == 124) || 
(treg[15:8] == 123 && freg[15:8] == 124) || 
(freg[15:8] == 124 && treg[15:8] == 125) || 
(treg[15:8] == 124 && freg[15:8] == 125) || 
(freg[15:8] == 125 && treg[15:8] == 126) || 
(treg[15:8] == 125 && freg[15:8] == 126) || 
(freg[15:8] == 126 && treg[15:8] == 127) || 
(treg[15:8] == 126 && freg[15:8] == 127) || 
(freg[15:8] == 127 && treg[15:8] == 128) || 
(treg[15:8] == 127 && freg[15:8] == 128) || 
(freg[15:8] == 128 && treg[15:8] == 129) || 
(treg[15:8] == 128 && freg[15:8] == 129) || 
(freg[15:8] == 129 && treg[15:8] == 130) || 
(treg[15:8] == 129 && freg[15:8] == 130) || 
(freg[15:8] == 130 && treg[15:8] == 131) || 
(treg[15:8] == 130 && freg[15:8] == 131) || 
(freg[15:8] == 131 && treg[15:8] == 132) || 
(treg[15:8] == 131 && freg[15:8] == 132) || 
(freg[15:8] == 132 && treg[15:8] == 133) || 
(treg[15:8] == 132 && freg[15:8] == 133) || 
(freg[15:8] == 133 && treg[15:8] == 134) || 
(treg[15:8] == 133 && freg[15:8] == 134) || 
(freg[15:8] == 134 && treg[15:8] == 135) || 
(treg[15:8] == 134 && freg[15:8] == 135) || 
(freg[15:8] == 135 && treg[15:8] == 136) || 
(treg[15:8] == 135 && freg[15:8] == 136) || 
(freg[15:8] == 136 && treg[15:8] == 137) || 
(treg[15:8] == 136 && freg[15:8] == 137) || 
(freg[15:8] == 137 && treg[15:8] == 138) || 
(treg[15:8] == 137 && freg[15:8] == 138) || 
(freg[15:8] == 138 && treg[15:8] == 139) || 
(treg[15:8] == 138 && freg[15:8] == 139) || 
(freg[15:8] == 139 && treg[15:8] == 140) || 
(treg[15:8] == 139 && freg[15:8] == 140) || 
(freg[15:8] == 140 && treg[15:8] == 141) || 
(treg[15:8] == 140 && freg[15:8] == 141) || 
(freg[15:8] == 141 && treg[15:8] == 142) || 
(treg[15:8] == 141 && freg[15:8] == 142) || 
(freg[15:8] == 142 && treg[15:8] == 143) || 
(treg[15:8] == 142 && freg[15:8] == 143) || 
(freg[15:8] == 143 && treg[15:8] == 144) || 
(treg[15:8] == 143 && freg[15:8] == 144) || 
(freg[15:8] == 144 && treg[15:8] == 145) || 
(treg[15:8] == 144 && freg[15:8] == 145) || 
(freg[15:8] == 145 && treg[15:8] == 146) || 
(treg[15:8] == 145 && freg[15:8] == 146) || 
(freg[15:8] == 146 && treg[15:8] == 147) || 
(treg[15:8] == 146 && freg[15:8] == 147) || 
(freg[15:8] == 147 && treg[15:8] == 148) || 
(treg[15:8] == 147 && freg[15:8] == 148) || 
(freg[15:8] == 148 && treg[15:8] == 149) || 
(treg[15:8] == 148 && freg[15:8] == 149) || 
(freg[15:8] == 149 && treg[15:8] == 150) || 
(treg[15:8] == 149 && freg[15:8] == 150) || 
(freg[15:8] == 150 && treg[15:8] == 151) || 
(treg[15:8] == 150 && freg[15:8] == 151) || 
(freg[15:8] == 151 && treg[15:8] == 152) || 
(treg[15:8] == 151 && freg[15:8] == 152) || 
(freg[15:8] == 152 && treg[15:8] == 153) || 
(treg[15:8] == 152 && freg[15:8] == 153) || 
(freg[15:8] == 153 && treg[15:8] == 154) || 
(treg[15:8] == 153 && freg[15:8] == 154) || 
(freg[15:8] == 154 && treg[15:8] == 155) || 
(treg[15:8] == 154 && freg[15:8] == 155) || 
(freg[15:8] == 155 && treg[15:8] == 156) || 
(treg[15:8] == 155 && freg[15:8] == 156) || 
(freg[15:8] == 156 && treg[15:8] == 157) || 
(treg[15:8] == 156 && freg[15:8] == 157) || 
(freg[15:8] == 157 && treg[15:8] == 158) || 
(treg[15:8] == 157 && freg[15:8] == 158) || 
(freg[15:8] == 158 && treg[15:8] == 159) || 
(treg[15:8] == 158 && freg[15:8] == 159) || 
(freg[15:8] == 159 && treg[15:8] == 160) || 
(treg[15:8] == 159 && freg[15:8] == 160) || 
(freg[15:8] == 160 && treg[15:8] == 161) || 
(treg[15:8] == 160 && freg[15:8] == 161) || 
(freg[15:8] == 161 && treg[15:8] == 162) || 
(treg[15:8] == 161 && freg[15:8] == 162) || 
(freg[15:8] == 162 && treg[15:8] == 163) || 
(treg[15:8] == 162 && freg[15:8] == 163) || 
(freg[15:8] == 163 && treg[15:8] == 164) || 
(treg[15:8] == 163 && freg[15:8] == 164) || 
(freg[15:8] == 164 && treg[15:8] == 165) || 
(treg[15:8] == 164 && freg[15:8] == 165) || 
(freg[15:8] == 165 && treg[15:8] == 166) || 
(treg[15:8] == 165 && freg[15:8] == 166) || 
(freg[15:8] == 166 && treg[15:8] == 167) || 
(treg[15:8] == 166 && freg[15:8] == 167) || 
(freg[15:8] == 167 && treg[15:8] == 168) || 
(treg[15:8] == 167 && freg[15:8] == 168) || 
(freg[15:8] == 168 && treg[15:8] == 169) || 
(treg[15:8] == 168 && freg[15:8] == 169) || 
(freg[15:8] == 169 && treg[15:8] == 170) || 
(treg[15:8] == 169 && freg[15:8] == 170) || 
(freg[15:8] == 170 && treg[15:8] == 171) || 
(treg[15:8] == 170 && freg[15:8] == 171) || 
(freg[15:8] == 171 && treg[15:8] == 172) || 
(treg[15:8] == 171 && freg[15:8] == 172) || 
(freg[15:8] == 172 && treg[15:8] == 173) || 
(treg[15:8] == 172 && freg[15:8] == 173) || 
(freg[15:8] == 173 && treg[15:8] == 174) || 
(treg[15:8] == 173 && freg[15:8] == 174) || 
(freg[15:8] == 174 && treg[15:8] == 175) || 
(treg[15:8] == 174 && freg[15:8] == 175) || 
(freg[15:8] == 175 && treg[15:8] == 176) || 
(treg[15:8] == 175 && freg[15:8] == 176) || 
(freg[15:8] == 176 && treg[15:8] == 177) || 
(treg[15:8] == 176 && freg[15:8] == 177) || 
(freg[15:8] == 177 && treg[15:8] == 178) || 
(treg[15:8] == 177 && freg[15:8] == 178) || 
(freg[15:8] == 178 && treg[15:8] == 179) || 
(treg[15:8] == 178 && freg[15:8] == 179) || 
(freg[15:8] == 179 && treg[15:8] == 180) || 
(treg[15:8] == 179 && freg[15:8] == 180) || 
(freg[15:8] == 180 && treg[15:8] == 181) || 
(treg[15:8] == 180 && freg[15:8] == 181) || 
(freg[15:8] == 181 && treg[15:8] == 182) || 
(treg[15:8] == 181 && freg[15:8] == 182) || 
(freg[15:8] == 182 && treg[15:8] == 183) || 
(treg[15:8] == 182 && freg[15:8] == 183) || 
(freg[15:8] == 183 && treg[15:8] == 184) || 
(treg[15:8] == 183 && freg[15:8] == 184) || 
(freg[15:8] == 184 && treg[15:8] == 185) || 
(treg[15:8] == 184 && freg[15:8] == 185) || 
(freg[15:8] == 185 && treg[15:8] == 186) || 
(treg[15:8] == 185 && freg[15:8] == 186) || 
(freg[15:8] == 186 && treg[15:8] == 187) || 
(treg[15:8] == 186 && freg[15:8] == 187) || 
(freg[15:8] == 187 && treg[15:8] == 188) || 
(treg[15:8] == 187 && freg[15:8] == 188) || 
(freg[15:8] == 188 && treg[15:8] == 189) || 
(treg[15:8] == 188 && freg[15:8] == 189) || 
(freg[15:8] == 189 && treg[15:8] == 190) || 
(treg[15:8] == 189 && freg[15:8] == 190) || 
(freg[15:8] == 190 && treg[15:8] == 191) || 
(treg[15:8] == 190 && freg[15:8] == 191) || 
(freg[15:8] == 191 && treg[15:8] == 192) || 
(treg[15:8] == 191 && freg[15:8] == 192) || 
(freg[15:8] == 192 && treg[15:8] == 193) || 
(treg[15:8] == 192 && freg[15:8] == 193) || 
(freg[15:8] == 193 && treg[15:8] == 194) || 
(treg[15:8] == 193 && freg[15:8] == 194) || 
(freg[15:8] == 194 && treg[15:8] == 195) || 
(treg[15:8] == 194 && freg[15:8] == 195) || 
(freg[15:8] == 195 && treg[15:8] == 196) || 
(treg[15:8] == 195 && freg[15:8] == 196) || 
(freg[15:8] == 196 && treg[15:8] == 197) || 
(treg[15:8] == 196 && freg[15:8] == 197) || 
(freg[15:8] == 197 && treg[15:8] == 198) || 
(treg[15:8] == 197 && freg[15:8] == 198) || 
(freg[15:8] == 198 && treg[15:8] == 199) || 
(treg[15:8] == 198 && freg[15:8] == 199) || 
(freg[15:8] == 199 && treg[15:8] == 200) || 
(treg[15:8] == 199 && freg[15:8] == 200) || 
(freg[15:8] == 200 && treg[15:8] == 201) || 
(treg[15:8] == 200 && freg[15:8] == 201) || 
(freg[15:8] == 201 && treg[15:8] == 202) || 
(treg[15:8] == 201 && freg[15:8] == 202) || 
(freg[15:8] == 202 && treg[15:8] == 203) || 
(treg[15:8] == 202 && freg[15:8] == 203) || 
(freg[15:8] == 203 && treg[15:8] == 204) || 
(treg[15:8] == 203 && freg[15:8] == 204) || 
(freg[15:8] == 204 && treg[15:8] == 205) || 
(treg[15:8] == 204 && freg[15:8] == 205) || 
(freg[15:8] == 205 && treg[15:8] == 206) || 
(treg[15:8] == 205 && freg[15:8] == 206) || 
(freg[15:8] == 206 && treg[15:8] == 207) || 
(treg[15:8] == 206 && freg[15:8] == 207) || 
(freg[15:8] == 207 && treg[15:8] == 208) || 
(treg[15:8] == 207 && freg[15:8] == 208) || 
(freg[15:8] == 208 && treg[15:8] == 209) || 
(treg[15:8] == 208 && freg[15:8] == 209) || 
(freg[15:8] == 209 && treg[15:8] == 210) || 
(treg[15:8] == 209 && freg[15:8] == 210) || 
(freg[15:8] == 210 && treg[15:8] == 211) || 
(treg[15:8] == 210 && freg[15:8] == 211) || 
(freg[15:8] == 211 && treg[15:8] == 212) || 
(treg[15:8] == 211 && freg[15:8] == 212) || 
(freg[15:8] == 212 && treg[15:8] == 213) || 
(treg[15:8] == 212 && freg[15:8] == 213) || 
(freg[15:8] == 213 && treg[15:8] == 214) || 
(treg[15:8] == 213 && freg[15:8] == 214) || 
(freg[15:8] == 214 && treg[15:8] == 215) || 
(treg[15:8] == 214 && freg[15:8] == 215) || 
(freg[15:8] == 215 && treg[15:8] == 216) || 
(treg[15:8] == 215 && freg[15:8] == 216) || 
(freg[15:8] == 216 && treg[15:8] == 217) || 
(treg[15:8] == 216 && freg[15:8] == 217) || 
(freg[15:8] == 217 && treg[15:8] == 218) || 
(treg[15:8] == 217 && freg[15:8] == 218) || 
(freg[15:8] == 218 && treg[15:8] == 219) || 
(treg[15:8] == 218 && freg[15:8] == 219) || 
(freg[15:8] == 219 && treg[15:8] == 220) || 
(treg[15:8] == 219 && freg[15:8] == 220) || 
(freg[15:8] == 220 && treg[15:8] == 221) || 
(treg[15:8] == 220 && freg[15:8] == 221) || 
(freg[15:8] == 221 && treg[15:8] == 222) || 
(treg[15:8] == 221 && freg[15:8] == 222) || 
(freg[15:8] == 222 && treg[15:8] == 223) || 
(treg[15:8] == 222 && freg[15:8] == 223) || 
(freg[15:8] == 223 && treg[15:8] == 224) || 
(treg[15:8] == 223 && freg[15:8] == 224) || 
(freg[15:8] == 224 && treg[15:8] == 225) || 
(treg[15:8] == 224 && freg[15:8] == 225) || 
(freg[15:8] == 225 && treg[15:8] == 226) || 
(treg[15:8] == 225 && freg[15:8] == 226) || 
(freg[15:8] == 226 && treg[15:8] == 227) || 
(treg[15:8] == 226 && freg[15:8] == 227) || 
(freg[15:8] == 227 && treg[15:8] == 228) || 
(treg[15:8] == 227 && freg[15:8] == 228) || 
(freg[15:8] == 228 && treg[15:8] == 229) || 
(treg[15:8] == 228 && freg[15:8] == 229) || 
(freg[15:8] == 229 && treg[15:8] == 230) || 
(treg[15:8] == 229 && freg[15:8] == 230) || 
(freg[15:8] == 230 && treg[15:8] == 231) || 
(treg[15:8] == 230 && freg[15:8] == 231) || 
(freg[15:8] == 231 && treg[15:8] == 232) || 
(treg[15:8] == 231 && freg[15:8] == 232) || 
(freg[15:8] == 232 && treg[15:8] == 233) || 
(treg[15:8] == 232 && freg[15:8] == 233) || 
(freg[15:8] == 233 && treg[15:8] == 234) || 
(treg[15:8] == 233 && freg[15:8] == 234) || 
(freg[15:8] == 234 && treg[15:8] == 235) || 
(treg[15:8] == 234 && freg[15:8] == 235) || 
(freg[15:8] == 235 && treg[15:8] == 236) || 
(treg[15:8] == 235 && freg[15:8] == 236) || 
(freg[15:8] == 236 && treg[15:8] == 237) || 
(treg[15:8] == 236 && freg[15:8] == 237) || 
(freg[15:8] == 237 && treg[15:8] == 238) || 
(treg[15:8] == 237 && freg[15:8] == 238) || 
(freg[15:8] == 238 && treg[15:8] == 239) || 
(treg[15:8] == 238 && freg[15:8] == 239) || 
(freg[15:8] == 239 && treg[15:8] == 240) || 
(treg[15:8] == 239 && freg[15:8] == 240) || 
(freg[15:8] == 240 && treg[15:8] == 241) || 
(treg[15:8] == 240 && freg[15:8] == 241) || 
(freg[15:8] == 241 && treg[15:8] == 242) || 
(treg[15:8] == 241 && freg[15:8] == 242) || 
(freg[15:8] == 242 && treg[15:8] == 243) || 
(treg[15:8] == 242 && freg[15:8] == 243) || 
(freg[15:8] == 243 && treg[15:8] == 244) || 
(treg[15:8] == 243 && freg[15:8] == 244) || 
(freg[15:8] == 244 && treg[15:8] == 245) || 
(treg[15:8] == 244 && freg[15:8] == 245) || 
(freg[15:8] == 245 && treg[15:8] == 246) || 
(treg[15:8] == 245 && freg[15:8] == 246) || 
(freg[15:8] == 246 && treg[15:8] == 247) || 
(treg[15:8] == 246 && freg[15:8] == 247) || 
(freg[15:8] == 247 && treg[15:8] == 248) || 
(treg[15:8] == 247 && freg[15:8] == 248) || 
(freg[15:8] == 248 && treg[15:8] == 249) || 
(treg[15:8] == 248 && freg[15:8] == 249) || 
(freg[15:8] == 249 && treg[15:8] == 250) || 
(treg[15:8] == 249 && freg[15:8] == 250) || 
(freg[15:8] == 250 && treg[15:8] == 251) || 
(treg[15:8] == 250 && freg[15:8] == 251) || 
(freg[15:8] == 251 && treg[15:8] == 252) || 
(treg[15:8] == 251 && freg[15:8] == 252) || 
(freg[15:8] == 252 && treg[15:8] == 253) || 
(treg[15:8] == 252 && freg[15:8] == 253) || 
(freg[15:8] == 253 && treg[15:8] == 254) || 
(treg[15:8] == 253 && freg[15:8] == 254) || 
(freg[15:8] == 254 && treg[15:8] == 255) || 
(treg[15:8] == 254 && freg[15:8] == 255) || 
(freg[15:8] == 255 && treg[15:8] == 256) || 
(treg[15:8] == 255 && freg[15:8] == 256) || 
(freg[15:8] == 256 && treg[15:8] == 257) || 
(treg[15:8] == 256 && freg[15:8] == 257) || 
(freg[15:8] == 257 && treg[15:8] == 258) || 
(treg[15:8] == 257 && freg[15:8] == 258) || 
(freg[15:8] == 258 && treg[15:8] == 259) || 
(treg[15:8] == 258 && freg[15:8] == 259) || 
(freg[15:8] == 259 && treg[15:8] == 260) || 
(treg[15:8] == 259 && freg[15:8] == 260) || 
(freg[15:8] == 260 && treg[15:8] == 261) || 
(treg[15:8] == 260 && freg[15:8] == 261) || 
(freg[15:8] == 261 && treg[15:8] == 262) || 
(treg[15:8] == 261 && freg[15:8] == 262) || 
(freg[15:8] == 262 && treg[15:8] == 263) || 
(treg[15:8] == 262 && freg[15:8] == 263) || 
(freg[15:8] == 253 && treg[15:8] == 254) || 
(treg[15:8] == 253 && freg[15:8] == 254) || 
(freg[15:8] == 254 && treg[15:8] == 255) || 
(treg[15:8] == 254 && freg[15:8] == 255)
 
)                        
                    ||    //sliding within rows
                   (treg[11:6] == freg[11:6] && ((freg[7:0] == 0 && treg[7:0] == 1) || 
(treg[7:0] == 0 && freg[7:0] == 1) || 
(freg[7:0] == 1 && treg[7:0] == 2) || 
(treg[7:0] == 1 && freg[7:0] == 2) || 
(freg[7:0] == 2 && treg[7:0] == 3) || 
(treg[7:0] == 2 && freg[7:0] == 3) || 
(freg[7:0] == 3 && treg[7:0] == 4) || 
(treg[7:0] == 3 && freg[7:0] == 4) || 
(freg[7:0] == 4 && treg[7:0] == 5) || 
(treg[7:0] == 4 && freg[7:0] == 5) || 
(freg[7:0] == 5 && treg[7:0] == 6) || 
(treg[7:0] == 5 && freg[7:0] == 6) || 
(freg[7:0] == 6 && treg[7:0] == 7) || 
(treg[7:0] == 6 && freg[7:0] == 7) || 
(freg[7:0] == 7 && treg[7:0] == 8) || 
(treg[7:0] == 7 && freg[7:0] == 8) || 
(freg[7:0] == 8 && treg[7:0] == 9) || 
(treg[7:0] == 8 && freg[7:0] == 9) || 
(freg[7:0] == 9 && treg[7:0] == 10) || 
(treg[7:0] == 9 && freg[7:0] == 10) || 
(freg[7:0] == 10 && treg[7:0] == 11) || 
(treg[7:0] == 10 && freg[7:0] == 11) || 
(freg[7:0] == 11 && treg[7:0] == 12) || 
(treg[7:0] == 11 && freg[7:0] == 12) || 
(freg[7:0] == 12 && treg[7:0] == 13) || 
(treg[7:0] == 12 && freg[7:0] == 13) || 
(freg[7:0] == 13 && treg[7:0] == 14) || 
(treg[7:0] == 13 && freg[7:0] == 14) || 
(freg[7:0] == 14 && treg[7:0] == 15) || 
(treg[7:0] == 14 && freg[7:0] == 15) || 
(freg[7:0] == 15 && treg[7:0] == 16) || 
(treg[7:0] == 15 && freg[7:0] == 16) || 
(freg[7:0] == 16 && treg[7:0] == 17) || 
(treg[7:0] == 16 && freg[7:0] == 17) || 
(freg[7:0] == 17 && treg[7:0] == 18) || 
(treg[7:0] == 17 && freg[7:0] == 18) || 
(freg[7:0] == 18 && treg[7:0] == 19) || 
(treg[7:0] == 18 && freg[7:0] == 19) || 
(freg[7:0] == 19 && treg[7:0] == 20) || 
(treg[7:0] == 19 && freg[7:0] == 20) || 
(freg[7:0] == 20 && treg[7:0] == 21) || 
(treg[7:0] == 20 && freg[7:0] == 21) || 
(freg[7:0] == 21 && treg[7:0] == 22) || 
(treg[7:0] == 21 && freg[7:0] == 22) || 
(freg[7:0] == 22 && treg[7:0] == 23) || 
(treg[7:0] == 22 && freg[7:0] == 23) || 
(freg[7:0] == 23 && treg[7:0] == 24) || 
(treg[7:0] == 23 && freg[7:0] == 24) || 
(freg[7:0] == 24 && treg[7:0] == 25) || 
(treg[7:0] == 24 && freg[7:0] == 25) || 
(freg[7:0] == 25 && treg[7:0] == 26) || 
(treg[7:0] == 25 && freg[7:0] == 26) || 
(freg[7:0] == 26 && treg[7:0] == 27) || 
(treg[7:0] == 26 && freg[7:0] == 27) || 
(freg[7:0] == 27 && treg[7:0] == 28) || 
(treg[7:0] == 27 && freg[7:0] == 28) || 
(freg[7:0] == 28 && treg[7:0] == 29) || 
(treg[7:0] == 28 && freg[7:0] == 29) || 
(freg[7:0] == 29 && treg[7:0] == 30) || 
(treg[7:0] == 29 && freg[7:0] == 30) || 
(freg[7:0] == 30 && treg[7:0] == 31) || 
(treg[7:0] == 30 && freg[7:0] == 31) || 
(freg[7:0] == 31 && treg[7:0] == 32) || 
(treg[7:0] == 31 && freg[7:0] == 32) || 
(freg[7:0] == 32 && treg[7:0] == 33) || 
(treg[7:0] == 32 && freg[7:0] == 33) || 
(freg[7:0] == 33 && treg[7:0] == 34) || 
(treg[7:0] == 33 && freg[7:0] == 34) || 
(freg[7:0] == 34 && treg[7:0] == 35) || 
(treg[7:0] == 34 && freg[7:0] == 35) || 
(freg[7:0] == 35 && treg[7:0] == 36) || 
(treg[7:0] == 35 && freg[7:0] == 36) || 
(freg[7:0] == 36 && treg[7:0] == 37) || 
(treg[7:0] == 36 && freg[7:0] == 37) || 
(freg[7:0] == 37 && treg[7:0] == 38) || 
(treg[7:0] == 37 && freg[7:0] == 38) || 
(freg[7:0] == 38 && treg[7:0] == 39) || 
(treg[7:0] == 38 && freg[7:0] == 39) || 
(freg[7:0] == 39 && treg[7:0] == 40) || 
(treg[7:0] == 39 && freg[7:0] == 40) || 
(freg[7:0] == 40 && treg[7:0] == 41) || 
(treg[7:0] == 40 && freg[7:0] == 41) || 
(freg[7:0] == 41 && treg[7:0] == 42) || 
(treg[7:0] == 41 && freg[7:0] == 42) || 
(freg[7:0] == 42 && treg[7:0] == 43) || 
(treg[7:0] == 42 && freg[7:0] == 43) || 
(freg[7:0] == 43 && treg[7:0] == 44) || 
(treg[7:0] == 43 && freg[7:0] == 44) || 
(freg[7:0] == 44 && treg[7:0] == 45) || 
(treg[7:0] == 44 && freg[7:0] == 45) || 
(freg[7:0] == 45 && treg[7:0] == 46) || 
(treg[7:0] == 45 && freg[7:0] == 46) || 
(freg[7:0] == 46 && treg[7:0] == 47) || 
(treg[7:0] == 46 && freg[7:0] == 47) || 
(freg[7:0] == 47 && treg[7:0] == 48) || 
(treg[7:0] == 47 && freg[7:0] == 48) || 
(freg[7:0] == 48 && treg[7:0] == 49) || 
(treg[7:0] == 48 && freg[7:0] == 49) || 
(freg[7:0] == 49 && treg[7:0] == 50) || 
(treg[7:0] == 49 && freg[7:0] == 50) || 
(freg[7:0] == 50 && treg[7:0] == 51) || 
(treg[7:0] == 50 && freg[7:0] == 51) || 
(freg[7:0] == 51 && treg[7:0] == 52) || 
(treg[7:0] == 51 && freg[7:0] == 52) || 
(freg[7:0] == 52 && treg[7:0] == 53) || 
(treg[7:0] == 52 && freg[7:0] == 53) || 
(freg[7:0] == 53 && treg[7:0] == 54) || 
(treg[7:0] == 53 && freg[7:0] == 54) || 
(freg[7:0] == 54 && treg[7:0] == 55) || 
(treg[7:0] == 54 && freg[7:0] == 55) || 
(freg[7:0] == 55 && treg[7:0] == 56) || 
(treg[7:0] == 55 && freg[7:0] == 56) || 
(freg[7:0] == 56 && treg[7:0] == 57) || 
(treg[7:0] == 56 && freg[7:0] == 57) || 
(freg[7:0] == 57 && treg[7:0] == 58) || 
(treg[7:0] == 57 && freg[7:0] == 58) || 
(freg[7:0] == 58 && treg[7:0] == 59) || 
(treg[7:0] == 58 && freg[7:0] == 59) || 
(freg[7:0] == 59 && treg[7:0] == 60) || 
(treg[7:0] == 59 && freg[7:0] == 60) || 
(freg[7:0] == 60 && treg[7:0] == 61) || 
(treg[7:0] == 60 && freg[7:0] == 61) || 
(freg[7:0] == 61 && treg[7:0] == 62) || 
(treg[7:0] == 61 && freg[7:0] == 62) || 
(freg[7:0] == 62 && treg[7:0] == 63) || 
(treg[7:0] == 62 && freg[7:0] == 63) || 
(freg[7:0] == 63 && treg[7:0] == 64) || 
(treg[7:0] == 63 && freg[7:0] == 64) || 
(freg[7:0] == 64 && treg[7:0] == 65) || 
(treg[7:0] == 64 && freg[7:0] == 65) || 
(freg[7:0] == 65 && treg[7:0] == 66) || 
(treg[7:0] == 65 && freg[7:0] == 66) || 
(freg[7:0] == 66 && treg[7:0] == 67) || 
(treg[7:0] == 66 && freg[7:0] == 67) || 
(freg[7:0] == 67 && treg[7:0] == 68) || 
(treg[7:0] == 67 && freg[7:0] == 68) || 
(freg[7:0] == 68 && treg[7:0] == 69) || 
(treg[7:0] == 68 && freg[7:0] == 69) || 
(freg[7:0] == 69 && treg[7:0] == 70) || 
(treg[7:0] == 69 && freg[7:0] == 70) || 
(freg[7:0] == 70 && treg[7:0] == 71) || 
(treg[7:0] == 70 && freg[7:0] == 71) || 
(freg[7:0] == 71 && treg[7:0] == 72) || 
(treg[7:0] == 71 && freg[7:0] == 72) || 
(freg[7:0] == 72 && treg[7:0] == 73) || 
(treg[7:0] == 72 && freg[7:0] == 73) || 
(freg[7:0] == 73 && treg[7:0] == 74) || 
(treg[7:0] == 73 && freg[7:0] == 74) || 
(freg[7:0] == 74 && treg[7:0] == 75) || 
(treg[7:0] == 74 && freg[7:0] == 75) || 
(freg[7:0] == 75 && treg[7:0] == 76) || 
(treg[7:0] == 75 && freg[7:0] == 76) || 
(freg[7:0] == 76 && treg[7:0] == 77) || 
(treg[7:0] == 76 && freg[7:0] == 77) || 
(freg[7:0] == 77 && treg[7:0] == 78) || 
(treg[7:0] == 77 && freg[7:0] == 78) || 
(freg[7:0] == 78 && treg[7:0] == 79) || 
(treg[7:0] == 78 && freg[7:0] == 79) || 
(freg[7:0] == 79 && treg[7:0] == 80) || 
(treg[7:0] == 79 && freg[7:0] == 80) || 
(freg[7:0] == 80 && treg[7:0] == 81) || 
(treg[7:0] == 80 && freg[7:0] == 81) || 
(freg[7:0] == 81 && treg[7:0] == 82) || 
(treg[7:0] == 81 && freg[7:0] == 82) || 
(freg[7:0] == 82 && treg[7:0] == 83) || 
(treg[7:0] == 82 && freg[7:0] == 83) || 
(freg[7:0] == 83 && treg[7:0] == 84) || 
(treg[7:0] == 83 && freg[7:0] == 84) || 
(freg[7:0] == 84 && treg[7:0] == 85) || 
(treg[7:0] == 84 && freg[7:0] == 85) || 
(freg[7:0] == 85 && treg[7:0] == 86) || 
(treg[7:0] == 85 && freg[7:0] == 86) || 
(freg[7:0] == 86 && treg[7:0] == 87) || 
(treg[7:0] == 86 && freg[7:0] == 87) || 
(freg[7:0] == 87 && treg[7:0] == 88) || 
(treg[7:0] == 87 && freg[7:0] == 88) || 
(freg[7:0] == 88 && treg[7:0] == 89) || 
(treg[7:0] == 88 && freg[7:0] == 89) || 
(freg[7:0] == 89 && treg[7:0] == 90) || 
(treg[7:0] == 89 && freg[7:0] == 90) || 
(freg[7:0] == 90 && treg[7:0] == 91) || 
(treg[7:0] == 90 && freg[7:0] == 91) || 
(freg[7:0] == 91 && treg[7:0] == 92) || 
(treg[7:0] == 91 && freg[7:0] == 92) || 
(freg[7:0] == 92 && treg[7:0] == 93) || 
(treg[7:0] == 92 && freg[7:0] == 93) || 
(freg[7:0] == 93 && treg[7:0] == 94) || 
(treg[7:0] == 93 && freg[7:0] == 94) || 
(freg[7:0] == 94 && treg[7:0] == 95) || 
(treg[7:0] == 94 && freg[7:0] == 95) || 
(freg[7:0] == 95 && treg[7:0] == 96) || 
(treg[7:0] == 95 && freg[7:0] == 96) || 
(freg[7:0] == 96 && treg[7:0] == 97) || 
(treg[7:0] == 96 && freg[7:0] == 97) || 
(freg[7:0] == 97 && treg[7:0] == 98) || 
(treg[7:0] == 97 && freg[7:0] == 98) || 
(freg[7:0] == 98 && treg[7:0] == 99) || 
(treg[7:0] == 98 && freg[7:0] == 99) || 
(freg[7:0] == 99 && treg[7:0] == 100) || 
(treg[7:0] == 99 && freg[7:0] == 100) || 
(freg[7:0] == 100 && treg[7:0] == 101) || 
(treg[7:0] == 100 && freg[7:0] == 101) || 
(freg[7:0] == 101 && treg[7:0] == 102) || 
(treg[7:0] == 101 && freg[7:0] == 102) || 
(freg[7:0] == 102 && treg[7:0] == 103) || 
(treg[7:0] == 102 && freg[7:0] == 103) || 
(freg[7:0] == 103 && treg[7:0] == 104) || 
(treg[7:0] == 103 && freg[7:0] == 104) || 
(freg[7:0] == 104 && treg[7:0] == 105) || 
(treg[7:0] == 104 && freg[7:0] == 105) || 
(freg[7:0] == 105 && treg[7:0] == 106) || 
(treg[7:0] == 105 && freg[7:0] == 106) || 
(freg[7:0] == 106 && treg[7:0] == 107) || 
(treg[7:0] == 106 && freg[7:0] == 107) || 
(freg[7:0] == 107 && treg[7:0] == 108) || 
(treg[7:0] == 107 && freg[7:0] == 108) || 
(freg[7:0] == 108 && treg[7:0] == 109) || 
(treg[7:0] == 108 && freg[7:0] == 109) || 
(freg[7:0] == 109 && treg[7:0] == 110) || 
(treg[7:0] == 109 && freg[7:0] == 110) || 
(freg[7:0] == 110 && treg[7:0] == 111) || 
(treg[7:0] == 110 && freg[7:0] == 111) || 
(freg[7:0] == 111 && treg[7:0] == 112) || 
(treg[7:0] == 111 && freg[7:0] == 112) || 
(freg[7:0] == 112 && treg[7:0] == 113) || 
(treg[7:0] == 112 && freg[7:0] == 113) || 
(freg[7:0] == 113 && treg[7:0] == 114) || 
(treg[7:0] == 113 && freg[7:0] == 114) || 
(freg[7:0] == 114 && treg[7:0] == 115) || 
(treg[7:0] == 114 && freg[7:0] == 115) || 
(freg[7:0] == 115 && treg[7:0] == 116) || 
(treg[7:0] == 115 && freg[7:0] == 116) || 
(freg[7:0] == 116 && treg[7:0] == 117) || 
(treg[7:0] == 116 && freg[7:0] == 117) || 
(freg[7:0] == 117 && treg[7:0] == 118) || 
(treg[7:0] == 117 && freg[7:0] == 118) || 
(freg[7:0] == 118 && treg[7:0] == 119) || 
(treg[7:0] == 118 && freg[7:0] == 119) || 
(freg[7:0] == 119 && treg[7:0] == 120) || 
(treg[7:0] == 119 && freg[7:0] == 120) || 
(freg[7:0] == 120 && treg[7:0] == 121) || 
(treg[7:0] == 120 && freg[7:0] == 121) || 
(freg[7:0] == 121 && treg[7:0] == 122) || 
(treg[7:0] == 121 && freg[7:0] == 122) || 
(freg[7:0] == 122 && treg[7:0] == 123) || 
(treg[7:0] == 122 && freg[7:0] == 123) || 
(freg[7:0] == 123 && treg[7:0] == 124) || 
(treg[7:0] == 123 && freg[7:0] == 124) || 
(freg[7:0] == 124 && treg[7:0] == 125) || 
(treg[7:0] == 124 && freg[7:0] == 125) || 
(freg[7:0] == 125 && treg[7:0] == 126) || 
(treg[7:0] == 125 && freg[7:0] == 126) || 
(freg[7:0] == 126 && treg[7:0] == 127) || 
(treg[7:0] == 126 && freg[7:0] == 127) || 
(freg[7:0] == 127 && treg[7:0] == 128) || 
(treg[7:0] == 127 && freg[7:0] == 128) || 
(freg[7:0] == 128 && treg[7:0] == 129) || 
(treg[7:0] == 128 && freg[7:0] == 129) || 
(freg[7:0] == 129 && treg[7:0] == 130) || 
(treg[7:0] == 129 && freg[7:0] == 130) || 
(freg[7:0] == 130 && treg[7:0] == 131) || 
(treg[7:0] == 130 && freg[7:0] == 131) || 
(freg[7:0] == 131 && treg[7:0] == 132) || 
(treg[7:0] == 131 && freg[7:0] == 132) || 
(freg[7:0] == 132 && treg[7:0] == 133) || 
(treg[7:0] == 132 && freg[7:0] == 133) || 
(freg[7:0] == 133 && treg[7:0] == 134) || 
(treg[7:0] == 133 && freg[7:0] == 134) || 
(freg[7:0] == 134 && treg[7:0] == 135) || 
(treg[7:0] == 134 && freg[7:0] == 135) || 
(freg[7:0] == 135 && treg[7:0] == 136) || 
(treg[7:0] == 135 && freg[7:0] == 136) || 
(freg[7:0] == 136 && treg[7:0] == 137) || 
(treg[7:0] == 136 && freg[7:0] == 137) || 
(freg[7:0] == 137 && treg[7:0] == 138) || 
(treg[7:0] == 137 && freg[7:0] == 138) || 
(freg[7:0] == 138 && treg[7:0] == 139) || 
(treg[7:0] == 138 && freg[7:0] == 139) || 
(freg[7:0] == 139 && treg[7:0] == 140) || 
(treg[7:0] == 139 && freg[7:0] == 140) || 
(freg[7:0] == 140 && treg[7:0] == 141) || 
(treg[7:0] == 140 && freg[7:0] == 141) || 
(freg[7:0] == 141 && treg[7:0] == 142) || 
(treg[7:0] == 141 && freg[7:0] == 142) || 
(freg[7:0] == 142 && treg[7:0] == 143) || 
(treg[7:0] == 142 && freg[7:0] == 143) || 
(freg[7:0] == 143 && treg[7:0] == 144) || 
(treg[7:0] == 143 && freg[7:0] == 144) || 
(freg[7:0] == 144 && treg[7:0] == 145) || 
(treg[7:0] == 144 && freg[7:0] == 145) || 
(freg[7:0] == 145 && treg[7:0] == 146) || 
(treg[7:0] == 145 && freg[7:0] == 146) || 
(freg[7:0] == 146 && treg[7:0] == 147) || 
(treg[7:0] == 146 && freg[7:0] == 147) || 
(freg[7:0] == 147 && treg[7:0] == 148) || 
(treg[7:0] == 147 && freg[7:0] == 148) || 
(freg[7:0] == 148 && treg[7:0] == 149) || 
(treg[7:0] == 148 && freg[7:0] == 149) || 
(freg[7:0] == 149 && treg[7:0] == 150) || 
(treg[7:0] == 149 && freg[7:0] == 150) || 
(freg[7:0] == 150 && treg[7:0] == 151) || 
(treg[7:0] == 150 && freg[7:0] == 151) || 
(freg[7:0] == 151 && treg[7:0] == 152) || 
(treg[7:0] == 151 && freg[7:0] == 152) || 
(freg[7:0] == 152 && treg[7:0] == 153) || 
(treg[7:0] == 152 && freg[7:0] == 153) || 
(freg[7:0] == 153 && treg[7:0] == 154) || 
(treg[7:0] == 153 && freg[7:0] == 154) || 
(freg[7:0] == 154 && treg[7:0] == 155) || 
(treg[7:0] == 154 && freg[7:0] == 155) || 
(freg[7:0] == 155 && treg[7:0] == 156) || 
(treg[7:0] == 155 && freg[7:0] == 156) || 
(freg[7:0] == 156 && treg[7:0] == 157) || 
(treg[7:0] == 156 && freg[7:0] == 157) || 
(freg[7:0] == 157 && treg[7:0] == 158) || 
(treg[7:0] == 157 && freg[7:0] == 158) || 
(freg[7:0] == 158 && treg[7:0] == 159) || 
(treg[7:0] == 158 && freg[7:0] == 159) || 
(freg[7:0] == 159 && treg[7:0] == 160) || 
(treg[7:0] == 159 && freg[7:0] == 160) || 
(freg[7:0] == 160 && treg[7:0] == 161) || 
(treg[7:0] == 160 && freg[7:0] == 161) || 
(freg[7:0] == 161 && treg[7:0] == 162) || 
(treg[7:0] == 161 && freg[7:0] == 162) || 
(freg[7:0] == 162 && treg[7:0] == 163) || 
(treg[7:0] == 162 && freg[7:0] == 163) || 
(freg[7:0] == 163 && treg[7:0] == 164) || 
(treg[7:0] == 163 && freg[7:0] == 164) || 
(freg[7:0] == 164 && treg[7:0] == 165) || 
(treg[7:0] == 164 && freg[7:0] == 165) || 
(freg[7:0] == 165 && treg[7:0] == 166) || 
(treg[7:0] == 165 && freg[7:0] == 166) || 
(freg[7:0] == 166 && treg[7:0] == 167) || 
(treg[7:0] == 166 && freg[7:0] == 167) || 
(freg[7:0] == 167 && treg[7:0] == 168) || 
(treg[7:0] == 167 && freg[7:0] == 168) || 
(freg[7:0] == 168 && treg[7:0] == 169) || 
(treg[7:0] == 168 && freg[7:0] == 169) || 
(freg[7:0] == 169 && treg[7:0] == 170) || 
(treg[7:0] == 169 && freg[7:0] == 170) || 
(freg[7:0] == 170 && treg[7:0] == 171) || 
(treg[7:0] == 170 && freg[7:0] == 171) || 
(freg[7:0] == 171 && treg[7:0] == 172) || 
(treg[7:0] == 171 && freg[7:0] == 172) || 
(freg[7:0] == 172 && treg[7:0] == 173) || 
(treg[7:0] == 172 && freg[7:0] == 173) || 
(freg[7:0] == 173 && treg[7:0] == 174) || 
(treg[7:0] == 173 && freg[7:0] == 174) || 
(freg[7:0] == 174 && treg[7:0] == 175) || 
(treg[7:0] == 174 && freg[7:0] == 175) || 
(freg[7:0] == 175 && treg[7:0] == 176) || 
(treg[7:0] == 175 && freg[7:0] == 176) || 
(freg[7:0] == 176 && treg[7:0] == 177) || 
(treg[7:0] == 176 && freg[7:0] == 177) || 
(freg[7:0] == 177 && treg[7:0] == 178) || 
(treg[7:0] == 177 && freg[7:0] == 178) || 
(freg[7:0] == 178 && treg[7:0] == 179) || 
(treg[7:0] == 178 && freg[7:0] == 179) || 
(freg[7:0] == 179 && treg[7:0] == 180) || 
(treg[7:0] == 179 && freg[7:0] == 180) || 
(freg[7:0] == 180 && treg[7:0] == 181) || 
(treg[7:0] == 180 && freg[7:0] == 181) || 
(freg[7:0] == 181 && treg[7:0] == 182) || 
(treg[7:0] == 181 && freg[7:0] == 182) || 
(freg[7:0] == 182 && treg[7:0] == 183) || 
(treg[7:0] == 182 && freg[7:0] == 183) || 
(freg[7:0] == 183 && treg[7:0] == 184) || 
(treg[7:0] == 183 && freg[7:0] == 184) || 
(freg[7:0] == 184 && treg[7:0] == 185) || 
(treg[7:0] == 184 && freg[7:0] == 185) || 
(freg[7:0] == 185 && treg[7:0] == 186) || 
(treg[7:0] == 185 && freg[7:0] == 186) || 
(freg[7:0] == 186 && treg[7:0] == 187) || 
(treg[7:0] == 186 && freg[7:0] == 187) || 
(freg[7:0] == 187 && treg[7:0] == 188) || 
(treg[7:0] == 187 && freg[7:0] == 188) || 
(freg[7:0] == 188 && treg[7:0] == 189) || 
(treg[7:0] == 188 && freg[7:0] == 189) || 
(freg[7:0] == 189 && treg[7:0] == 190) || 
(treg[7:0] == 189 && freg[7:0] == 190) || 
(freg[7:0] == 190 && treg[7:0] == 191) || 
(treg[7:0] == 190 && freg[7:0] == 191) || 
(freg[7:0] == 191 && treg[7:0] == 192) || 
(treg[7:0] == 191 && freg[7:0] == 192) || 
(freg[7:0] == 192 && treg[7:0] == 193) || 
(treg[7:0] == 192 && freg[7:0] == 193) || 
(freg[7:0] == 193 && treg[7:0] == 194) || 
(treg[7:0] == 193 && freg[7:0] == 194) || 
(freg[7:0] == 194 && treg[7:0] == 195) || 
(treg[7:0] == 194 && freg[7:0] == 195) || 
(freg[7:0] == 195 && treg[7:0] == 196) || 
(treg[7:0] == 195 && freg[7:0] == 196) || 
(freg[7:0] == 196 && treg[7:0] == 197) || 
(treg[7:0] == 196 && freg[7:0] == 197) || 
(freg[7:0] == 197 && treg[7:0] == 198) || 
(treg[7:0] == 197 && freg[7:0] == 198) || 
(freg[7:0] == 198 && treg[7:0] == 199) || 
(treg[7:0] == 198 && freg[7:0] == 199) || 
(freg[7:0] == 199 && treg[7:0] == 200) || 
(treg[7:0] == 199 && freg[7:0] == 200) || 
(freg[7:0] == 200 && treg[7:0] == 201) || 
(treg[7:0] == 200 && freg[7:0] == 201) || 
(freg[7:0] == 201 && treg[7:0] == 202) || 
(treg[7:0] == 201 && freg[7:0] == 202) || 
(freg[7:0] == 202 && treg[7:0] == 203) || 
(treg[7:0] == 202 && freg[7:0] == 203) || 
(freg[7:0] == 203 && treg[7:0] == 204) || 
(treg[7:0] == 203 && freg[7:0] == 204) || 
(freg[7:0] == 204 && treg[7:0] == 205) || 
(treg[7:0] == 204 && freg[7:0] == 205) || 
(freg[7:0] == 205 && treg[7:0] == 206) || 
(treg[7:0] == 205 && freg[7:0] == 206) || 
(freg[7:0] == 206 && treg[7:0] == 207) || 
(treg[7:0] == 206 && freg[7:0] == 207) || 
(freg[7:0] == 207 && treg[7:0] == 208) || 
(treg[7:0] == 207 && freg[7:0] == 208) || 
(freg[7:0] == 208 && treg[7:0] == 209) || 
(treg[7:0] == 208 && freg[7:0] == 209) || 
(freg[7:0] == 209 && treg[7:0] == 210) || 
(treg[7:0] == 209 && freg[7:0] == 210) || 
(freg[7:0] == 210 && treg[7:0] == 211) || 
(treg[7:0] == 210 && freg[7:0] == 211) || 
(freg[7:0] == 211 && treg[7:0] == 212) || 
(treg[7:0] == 211 && freg[7:0] == 212) || 
(freg[7:0] == 212 && treg[7:0] == 213) || 
(treg[7:0] == 212 && freg[7:0] == 213) || 
(freg[7:0] == 213 && treg[7:0] == 214) || 
(treg[7:0] == 213 && freg[7:0] == 214) || 
(freg[7:0] == 214 && treg[7:0] == 215) || 
(treg[7:0] == 214 && freg[7:0] == 215) || 
(freg[7:0] == 215 && treg[7:0] == 216) || 
(treg[7:0] == 215 && freg[7:0] == 216) || 
(freg[7:0] == 216 && treg[7:0] == 217) || 
(treg[7:0] == 216 && freg[7:0] == 217) || 
(freg[7:0] == 217 && treg[7:0] == 218) || 
(treg[7:0] == 217 && freg[7:0] == 218) || 
(freg[7:0] == 218 && treg[7:0] == 219) || 
(treg[7:0] == 218 && freg[7:0] == 219) || 
(freg[7:0] == 219 && treg[7:0] == 220) || 
(treg[7:0] == 219 && freg[7:0] == 220) || 
(freg[7:0] == 220 && treg[7:0] == 221) || 
(treg[7:0] == 220 && freg[7:0] == 221) || 
(freg[7:0] == 221 && treg[7:0] == 222) || 
(treg[7:0] == 221 && freg[7:0] == 222) || 
(freg[7:0] == 222 && treg[7:0] == 223) || 
(treg[7:0] == 222 && freg[7:0] == 223) || 
(freg[7:0] == 223 && treg[7:0] == 224) || 
(treg[7:0] == 223 && freg[7:0] == 224) || 
(freg[7:0] == 224 && treg[7:0] == 225) || 
(treg[7:0] == 224 && freg[7:0] == 225) || 
(freg[7:0] == 225 && treg[7:0] == 226) || 
(treg[7:0] == 225 && freg[7:0] == 226) || 
(freg[7:0] == 226 && treg[7:0] == 227) || 
(treg[7:0] == 226 && freg[7:0] == 227) || 
(freg[7:0] == 227 && treg[7:0] == 228) || 
(treg[7:0] == 227 && freg[7:0] == 228) || 
(freg[7:0] == 228 && treg[7:0] == 229) || 
(treg[7:0] == 228 && freg[7:0] == 229) || 
(freg[7:0] == 229 && treg[7:0] == 230) || 
(treg[7:0] == 229 && freg[7:0] == 230) || 
(freg[7:0] == 230 && treg[7:0] == 231) || 
(treg[7:0] == 230 && freg[7:0] == 231) || 
(freg[7:0] == 231 && treg[7:0] == 232) || 
(treg[7:0] == 231 && freg[7:0] == 232) || 
(freg[7:0] == 232 && treg[7:0] == 233) || 
(treg[7:0] == 232 && freg[7:0] == 233) || 
(freg[7:0] == 233 && treg[7:0] == 234) || 
(treg[7:0] == 233 && freg[7:0] == 234) || 
(freg[7:0] == 234 && treg[7:0] == 235) || 
(treg[7:0] == 234 && freg[7:0] == 235) || 
(freg[7:0] == 235 && treg[7:0] == 236) || 
(treg[7:0] == 235 && freg[7:0] == 236) || 
(freg[7:0] == 236 && treg[7:0] == 237) || 
(treg[7:0] == 236 && freg[7:0] == 237) || 
(freg[7:0] == 237 && treg[7:0] == 238) || 
(treg[7:0] == 237 && freg[7:0] == 238) || 
(freg[7:0] == 238 && treg[7:0] == 239) || 
(treg[7:0] == 238 && freg[7:0] == 239) || 
(freg[7:0] == 239 && treg[7:0] == 240) || 
(treg[7:0] == 239 && freg[7:0] == 240) || 
(freg[7:0] == 240 && treg[7:0] == 241) || 
(treg[7:0] == 240 && freg[7:0] == 241) || 
(freg[7:0] == 241 && treg[7:0] == 242) || 
(treg[7:0] == 241 && freg[7:0] == 242) || 
(freg[7:0] == 242 && treg[7:0] == 243) || 
(treg[7:0] == 242 && freg[7:0] == 243) || 
(freg[7:0] == 243 && treg[7:0] == 244) || 
(treg[7:0] == 243 && freg[7:0] == 244) || 
(freg[7:0] == 244 && treg[7:0] == 245) || 
(treg[7:0] == 244 && freg[7:0] == 245) || 
(freg[7:0] == 245 && treg[7:0] == 246) || 
(treg[7:0] == 245 && freg[7:0] == 246) || 
(freg[7:0] == 246 && treg[7:0] == 247) || 
(treg[7:0] == 246 && freg[7:0] == 247) || 
(freg[7:0] == 247 && treg[7:0] == 248) || 
(treg[7:0] == 247 && freg[7:0] == 248) || 
(freg[7:0] == 248 && treg[7:0] == 249) || 
(treg[7:0] == 248 && freg[7:0] == 249) || 
(freg[7:0] == 249 && treg[7:0] == 250) || 
(treg[7:0] == 249 && freg[7:0] == 250) || 
(freg[7:0] == 250 && treg[7:0] == 251) || 
(treg[7:0] == 250 && freg[7:0] == 251) || 
(freg[7:0] == 251 && treg[7:0] == 252) || 
(treg[7:0] == 251 && freg[7:0] == 252) || 
(freg[7:0] == 252 && treg[7:0] == 253) || 
(treg[7:0] == 252 && freg[7:0] == 253) || 
(freg[7:0] == 253 && treg[7:0] == 254) || 
(treg[7:0] == 253 && freg[7:0] == 254) || 
(freg[7:0] == 254 && treg[7:0] == 255) || 
(treg[7:0] == 254 && freg[7:0] == 255)

 )))
                     );
    assign parity = 
	   (((b[0] & 5) == 1) | ((b[0] & 5) == 4)) ^
	   (((b[1] & 5) == 0) | ((b[1] & 5) == 5)) ^
	   (((b[2] & 5) == 1) | ((b[2] & 5) == 4)) ^
	   (((b[3] & 5) == 0) | ((b[3] & 5) == 5)) ^
	   (((b[4] & 5) == 1) | ((b[4] & 5) == 4)) ^
	   (((b[5] & 5) == 0) | ((b[5] & 5) == 5)) ^
	   (((b[6] & 5) == 1) | ((b[6] & 5) == 4)) ^
	   (((b[7] & 5) == 0) | ((b[7] & 5) == 5));
 
    always @(posedge clock) begin
	freg <= from;
	treg <= to;
    end

    always @(posedge clock) begin
	if (valid) begin
	    b[treg] <= b[freg];
	    b[freg] <= 0;
	end
    end


logic [65535:0] match_bits;
genvar i;
    generate
        for (i = 0; i < 65536; i = i + 1) begin : gen_check
            always_comb match_bits[i] = (b[i] == i);
        end
    endgenerate

wire prop = ($countones(match_bits) == 65536);
assert property (@(posedge clock) !prop);

/*invariant property
!(b<*0*>[2:0]=0 * b<*1*>[2:0]=1 * b<*2*>[2:0]=2 * b<*3*>[2:0]=3 *
  b<*4*>[2:0]=4 * b<*5*>[2:0]=5 * b<*6*>[2:0]=6 * b<*7*>[2:0]=7);*/ 



endmodule //sliding_board
