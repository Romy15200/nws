/*
*
*	Taken from VIS Benchmarks <ftp://vlsi.colorado.edu/pub/vis/vis-verilog-models-1.3.tar.gz>
*	Modified by Ahmed Irfan <irfan@fbk.eu>
*
*/
//Author: Fabio Somenzi <Fabio@Colorado.EDU>
// Slider puzzle with N rows and N columns.             +-------+----+----+----+-----+-----+
//                                                      |  0    |  1 |  2 |  3 |.....| N-1 |
// The entries of the matrix are numbered thus:         +-------+----+----+----+-----+-----+
//                                                      |  N    | N+1| N+2| N+3|.....| 2N-1|
//                                                      +-------+----+----+----+-----+-----+  
//                                                      |.......|....|....|....|.....|.....|          
//                                                      +-------+----+----+----+-----+-----+
//                                                      |(N-1)*N|....|....|....|.....|N^2-1|
//                                                      +-------+----+----+----+-----+-----+
module slidingBoard(clock,from,to);
    input       clock;
    input [15:0] from;
    input [15:0] to;

    reg [15:0] 	b[0:65536];
    reg [15:0] 	freg, treg;
    wire 	valid, parity;

    initial begin
        for (i=0; i < 65536; i = i+1) begin
          b[i] = 65535-i;
	end
        treg = 0;
	freg = 0;
    end 

    assign valid = (b[treg] == 16'b0) &&
                    ( //sliding between rows
		   (treg[5:0] == freg[5:0] && ((freg[15:8] == 0 && treg[15:8] == 1) || 
(treg[15:8] == 0 && freg[15:8] == 1) || 
(freg[15:8] == 1 && treg[15:8] == 2) || 
(treg[15:8] == 1 && freg[15:8] == 2) || 
(freg[15:8] == 2 && treg[15:8] == 3) || 
(treg[15:8] == 2 && freg[15:8] == 3) || 
(freg[15:8] == 3 && treg[15:8] == 4) || 
(treg[15:8] == 3 && freg[15:8] == 4) || 
(freg[15:8] == 4 && treg[15:8] == 5) || 
(treg[15:8] == 4 && freg[15:8] == 5) || 
(freg[15:8] == 5 && treg[15:8] == 6) || 
(treg[15:8] == 5 && freg[15:8] == 6) || 
(freg[15:8] == 6 && treg[15:8] == 7) || 
(treg[15:8] == 6 && freg[15:8] == 7) || 
(freg[15:8] == 7 && treg[15:8] == 8) || 
(treg[15:8] == 7 && freg[15:8] == 8) || 
(freg[15:8] == 8 && treg[15:8] == 9) || 
(treg[15:8] == 8 && freg[15:8] == 9) || 
(freg[15:8] == 9 && treg[15:8] == 10) || 
(treg[15:8] == 9 && freg[15:8] == 10) || 
(freg[15:8] == 10 && treg[15:8] == 11) || 
(treg[15:8] == 10 && freg[15:8] == 11) || 
(freg[15:8] == 11 && treg[15:8] == 12) || 
(treg[15:8] == 11 && freg[15:8] == 12) || 
(freg[15:8] == 12 && treg[15:8] == 13) || 
(treg[15:8] == 12 && freg[15:8] == 13) || 
(freg[15:8] == 13 && treg[15:8] == 14) || 
(treg[15:8] == 13 && freg[15:8] == 14) || 
(freg[15:8] == 14 && treg[15:8] == 15) || 
(treg[15:8] == 14 && freg[15:8] == 15) || 
(freg[15:8] == 15 && treg[15:8] == 16) || 
(treg[15:8] == 15 && freg[15:8] == 16) || 
(freg[15:8] == 16 && treg[15:8] == 17) || 
(treg[15:8] == 16 && freg[15:8] == 17) || 
(freg[15:8] == 17 && treg[15:8] == 18) || 
(treg[15:8] == 17 && freg[15:8] == 18) || 
(freg[15:8] == 18 && treg[15:8] == 19) || 
(treg[15:8] == 18 && freg[15:8] == 19) || 
(freg[15:8] == 19 && treg[15:8] == 20) || 
(treg[15:8] == 19 && freg[15:8] == 20) || 
(freg[15:8] == 20 && treg[15:8] == 21) || 
(treg[15:8] == 20 && freg[15:8] == 21) || 
(freg[15:8] == 21 && treg[15:8] == 22) || 
(treg[15:8] == 21 && freg[15:8] == 22) || 
(freg[15:8] == 22 && treg[15:8] == 23) || 
(treg[15:8] == 22 && freg[15:8] == 23) || 
(freg[15:8] == 23 && treg[15:8] == 24) || 
(treg[15:8] == 23 && freg[15:8] == 24) || 
(freg[15:8] == 24 && treg[15:8] == 25) || 
(treg[15:8] == 24 && freg[15:8] == 25) || 
(freg[15:8] == 25 && treg[15:8] == 26) || 
(treg[15:8] == 25 && freg[15:8] == 26) || 
(freg[15:8] == 26 && treg[15:8] == 27) || 
(treg[15:8] == 26 && freg[15:8] == 27) || 
(freg[15:8] == 27 && treg[15:8] == 28) || 
(treg[15:8] == 27 && freg[15:8] == 28) || 
(freg[15:8] == 28 && treg[15:8] == 29) || 
(treg[15:8] == 28 && freg[15:8] == 29) || 
(freg[15:8] == 29 && treg[15:8] == 30) || 
(treg[15:8] == 29 && freg[15:8] == 30) || 
(freg[15:8] == 30 && treg[15:8] == 31) || 
(treg[15:8] == 30 && freg[15:8] == 31) || 
(freg[15:8] == 31 && treg[15:8] == 32) || 
(treg[15:8] == 31 && freg[15:8] == 32) || 
(freg[15:8] == 32 && treg[15:8] == 33) || 
(treg[15:8] == 32 && freg[15:8] == 33) || 
(freg[15:8] == 33 && treg[15:8] == 34) || 
(treg[15:8] == 33 && freg[15:8] == 34) || 
(freg[15:8] == 34 && treg[15:8] == 35) || 
(treg[15:8] == 34 && freg[15:8] == 35) || 
(freg[15:8] == 35 && treg[15:8] == 36) || 
(treg[15:8] == 35 && freg[15:8] == 36) || 
(freg[15:8] == 36 && treg[15:8] == 37) || 
(treg[15:8] == 36 && freg[15:8] == 37) || 
(freg[15:8] == 37 && treg[15:8] == 38) || 
(treg[15:8] == 37 && freg[15:8] == 38) || 
(freg[15:8] == 38 && treg[15:8] == 39) || 
(treg[15:8] == 38 && freg[15:8] == 39) || 
(freg[15:8] == 39 && treg[15:8] == 40) || 
(treg[15:8] == 39 && freg[15:8] == 40) || 
(freg[15:8] == 40 && treg[15:8] == 41) || 
(treg[15:8] == 40 && freg[15:8] == 41) || 
(freg[15:8] == 41 && treg[15:8] == 42) || 
(treg[15:8] == 41 && freg[15:8] == 42) || 
(freg[15:8] == 42 && treg[15:8] == 43) || 
(treg[15:8] == 42 && freg[15:8] == 43) || 
(freg[15:8] == 43 && treg[15:8] == 44) || 
(treg[15:8] == 43 && freg[15:8] == 44) || 
(freg[15:8] == 44 && treg[15:8] == 45) || 
(treg[15:8] == 44 && freg[15:8] == 45) || 
(freg[15:8] == 45 && treg[15:8] == 46) || 
(treg[15:8] == 45 && freg[15:8] == 46) || 
(freg[15:8] == 46 && treg[15:8] == 47) || 
(treg[15:8] == 46 && freg[15:8] == 47) || 
(freg[15:8] == 47 && treg[15:8] == 48) || 
(treg[15:8] == 47 && freg[15:8] == 48) || 
(freg[15:8] == 48 && treg[15:8] == 49) || 
(treg[15:8] == 48 && freg[15:8] == 49) || 
(freg[15:8] == 49 && treg[15:8] == 50) || 
(treg[15:8] == 49 && freg[15:8] == 50) || 
(freg[15:8] == 50 && treg[15:8] == 51) || 
(treg[15:8] == 50 && freg[15:8] == 51) || 
(freg[15:8] == 51 && treg[15:8] == 52) || 
(treg[15:8] == 51 && freg[15:8] == 52) || 
(freg[15:8] == 52 && treg[15:8] == 53) || 
(treg[15:8] == 52 && freg[15:8] == 53) || 
(freg[15:8] == 53 && treg[15:8] == 54) || 
(treg[15:8] == 53 && freg[15:8] == 54) || 
(freg[15:8] == 54 && treg[15:8] == 55) || 
(treg[15:8] == 54 && freg[15:8] == 55) || 
(freg[15:8] == 55 && treg[15:8] == 56) || 
(treg[15:8] == 55 && freg[15:8] == 56) || 
(freg[15:8] == 56 && treg[15:8] == 57) || 
(treg[15:8] == 56 && freg[15:8] == 57) || 
(freg[15:8] == 57 && treg[15:8] == 58) || 
(treg[15:8] == 57 && freg[15:8] == 58) || 
(freg[15:8] == 58 && treg[15:8] == 59) || 
(treg[15:8] == 58 && freg[15:8] == 59) || 
(freg[15:8] == 59 && treg[15:8] == 60) || 
(treg[15:8] == 59 && freg[15:8] == 60) || 
(freg[15:8] == 60 && treg[15:8] == 61) || 
(treg[15:8] == 60 && freg[15:8] == 61) || 
(freg[15:8] == 61 && treg[15:8] == 62) || 
(treg[15:8] == 61 && freg[15:8] == 62) || 
(freg[15:8] == 62 && treg[15:8] == 63) || 
(treg[15:8] == 62 && freg[15:8] == 63) || 
(freg[15:8] == 63 && treg[15:8] == 64) || 
(treg[15:8] == 63 && freg[15:8] == 64) || 
(freg[15:8] == 64 && treg[15:8] == 65) || 
(treg[15:8] == 64 && freg[15:8] == 65) || 
(freg[15:8] == 65 && treg[15:8] == 66) || 
(treg[15:8] == 65 && freg[15:8] == 66) || 
(freg[15:8] == 66 && treg[15:8] == 67) || 
(treg[15:8] == 66 && freg[15:8] == 67) || 
(freg[15:8] == 67 && treg[15:8] == 68) || 
(treg[15:8] == 67 && freg[15:8] == 68) || 
(freg[15:8] == 68 && treg[15:8] == 69) || 
(treg[15:8] == 68 && freg[15:8] == 69) || 
(freg[15:8] == 69 && treg[15:8] == 70) || 
(treg[15:8] == 69 && freg[15:8] == 70) || 
(freg[15:8] == 70 && treg[15:8] == 71) || 
(treg[15:8] == 70 && freg[15:8] == 71) || 
(freg[15:8] == 71 && treg[15:8] == 72) || 
(treg[15:8] == 71 && freg[15:8] == 72) || 
(freg[15:8] == 72 && treg[15:8] == 73) || 
(treg[15:8] == 72 && freg[15:8] == 73) || 
(freg[15:8] == 73 && treg[15:8] == 74) || 
(treg[15:8] == 73 && freg[15:8] == 74) || 
(freg[15:8] == 74 && treg[15:8] == 75) || 
(treg[15:8] == 74 && freg[15:8] == 75) || 
(freg[15:8] == 75 && treg[15:8] == 76) || 
(treg[15:8] == 75 && freg[15:8] == 76) || 
(freg[15:8] == 76 && treg[15:8] == 77) || 
(treg[15:8] == 76 && freg[15:8] == 77) || 
(freg[15:8] == 77 && treg[15:8] == 78) || 
(treg[15:8] == 77 && freg[15:8] == 78) || 
(freg[15:8] == 78 && treg[15:8] == 79) || 
(treg[15:8] == 78 && freg[15:8] == 79) || 
(freg[15:8] == 79 && treg[15:8] == 80) || 
(treg[15:8] == 79 && freg[15:8] == 80) || 
(freg[15:8] == 80 && treg[15:8] == 81) || 
(treg[15:8] == 80 && freg[15:8] == 81) || 
(freg[15:8] == 81 && treg[15:8] == 82) || 
(treg[15:8] == 81 && freg[15:8] == 82) || 
(freg[15:8] == 82 && treg[15:8] == 83) || 
(treg[15:8] == 82 && freg[15:8] == 83) || 
(freg[15:8] == 83 && treg[15:8] == 84) || 
(treg[15:8] == 83 && freg[15:8] == 84) || 
(freg[15:8] == 84 && treg[15:8] == 85) || 
(treg[15:8] == 84 && freg[15:8] == 85) || 
(freg[15:8] == 85 && treg[15:8] == 86) || 
(treg[15:8] == 85 && freg[15:8] == 86) || 
(freg[15:8] == 86 && treg[15:8] == 87) || 
(treg[15:8] == 86 && freg[15:8] == 87) || 
(freg[15:8] == 87 && treg[15:8] == 88) || 
(treg[15:8] == 87 && freg[15:8] == 88) || 
(freg[15:8] == 88 && treg[15:8] == 89) || 
(treg[15:8] == 88 && freg[15:8] == 89) || 
(freg[15:8] == 89 && treg[15:8] == 90) || 
(treg[15:8] == 89 && freg[15:8] == 90) || 
(freg[15:8] == 90 && treg[15:8] == 91) || 
(treg[15:8] == 90 && freg[15:8] == 91) || 
(freg[15:8] == 91 && treg[15:8] == 92) || 
(treg[15:8] == 91 && freg[15:8] == 92) || 
(freg[15:8] == 92 && treg[15:8] == 93) || 
(treg[15:8] == 92 && freg[15:8] == 93) || 
(freg[15:8] == 93 && treg[15:8] == 94) || 
(treg[15:8] == 93 && freg[15:8] == 94) || 
(freg[15:8] == 94 && treg[15:8] == 95) || 
(treg[15:8] == 94 && freg[15:8] == 95) || 
(freg[15:8] == 95 && treg[15:8] == 96) || 
(treg[15:8] == 95 && freg[15:8] == 96) || 
(freg[15:8] == 96 && treg[15:8] == 97) || 
(treg[15:8] == 96 && freg[15:8] == 97) || 
(freg[15:8] == 97 && treg[15:8] == 98) || 
(treg[15:8] == 97 && freg[15:8] == 98) || 
(freg[15:8] == 98 && treg[15:8] == 99) || 
(treg[15:8] == 98 && freg[15:8] == 99) || 
(freg[15:8] == 99 && treg[15:8] == 100) || 
(treg[15:8] == 99 && freg[15:8] == 100) || 
(freg[15:8] == 100 && treg[15:8] == 101) || 
(treg[15:8] == 100 && freg[15:8] == 101) || 
(freg[15:8] == 101 && treg[15:8] == 102) || 
(treg[15:8] == 101 && freg[15:8] == 102) || 
(freg[15:8] == 102 && treg[15:8] == 103) || 
(treg[15:8] == 102 && freg[15:8] == 103) || 
(freg[15:8] == 103 && treg[15:8] == 104) || 
(treg[15:8] == 103 && freg[15:8] == 104) || 
(freg[15:8] == 104 && treg[15:8] == 105) || 
(treg[15:8] == 104 && freg[15:8] == 105) || 
(freg[15:8] == 105 && treg[15:8] == 106) || 
(treg[15:8] == 105 && freg[15:8] == 106) || 
(freg[15:8] == 106 && treg[15:8] == 107) || 
(treg[15:8] == 106 && freg[15:8] == 107) || 
(freg[15:8] == 107 && treg[15:8] == 108) || 
(treg[15:8] == 107 && freg[15:8] == 108) || 
(freg[15:8] == 108 && treg[15:8] == 109) || 
(treg[15:8] == 108 && freg[15:8] == 109) || 
(freg[15:8] == 109 && treg[15:8] == 110) || 
(treg[15:8] == 109 && freg[15:8] == 110) || 
(freg[15:8] == 110 && treg[15:8] == 111) || 
(treg[15:8] == 110 && freg[15:8] == 111) || 
(freg[15:8] == 111 && treg[15:8] == 112) || 
(treg[15:8] == 111 && freg[15:8] == 112) || 
(freg[15:8] == 112 && treg[15:8] == 113) || 
(treg[15:8] == 112 && freg[15:8] == 113) || 
(freg[15:8] == 113 && treg[15:8] == 114) || 
(treg[15:8] == 113 && freg[15:8] == 114) || 
(freg[15:8] == 114 && treg[15:8] == 115) || 
(treg[15:8] == 114 && freg[15:8] == 115) || 
(freg[15:8] == 115 && treg[15:8] == 116) || 
(treg[15:8] == 115 && freg[15:8] == 116) || 
(freg[15:8] == 116 && treg[15:8] == 117) || 
(treg[15:8] == 116 && freg[15:8] == 117) || 
(freg[15:8] == 117 && treg[15:8] == 118) || 
(treg[15:8] == 117 && freg[15:8] == 118) || 
(freg[15:8] == 118 && treg[15:8] == 119) || 
(treg[15:8] == 118 && freg[15:8] == 119) || 
(freg[15:8] == 119 && treg[15:8] == 120) || 
(treg[15:8] == 119 && freg[15:8] == 120) || 
(freg[15:8] == 120 && treg[15:8] == 121) || 
(treg[15:8] == 120 && freg[15:8] == 121) || 
(freg[15:8] == 121 && treg[15:8] == 122) || 
(treg[15:8] == 121 && freg[15:8] == 122) || 
(freg[15:8] == 122 && treg[15:8] == 123) || 
(treg[15:8] == 122 && freg[15:8] == 123) || 
(freg[15:8] == 123 && treg[15:8] == 124) || 
(treg[15:8] == 123 && freg[15:8] == 124) || 
(freg[15:8] == 124 && treg[15:8] == 125) || 
(treg[15:8] == 124 && freg[15:8] == 125) || 
(freg[15:8] == 125 && treg[15:8] == 126) || 
(treg[15:8] == 125 && freg[15:8] == 126) || 
(freg[15:8] == 126 && treg[15:8] == 127) || 
(treg[15:8] == 126 && freg[15:8] == 127) || 
(freg[15:8] == 127 && treg[15:8] == 128) || 
(treg[15:8] == 127 && freg[15:8] == 128) || 
(freg[15:8] == 128 && treg[15:8] == 129) || 
(treg[15:8] == 128 && freg[15:8] == 129) || 
(freg[15:8] == 129 && treg[15:8] == 130) || 
(treg[15:8] == 129 && freg[15:8] == 130) || 
(freg[15:8] == 130 && treg[15:8] == 131) || 
(treg[15:8] == 130 && freg[15:8] == 131) || 
(freg[15:8] == 131 && treg[15:8] == 132) || 
(treg[15:8] == 131 && freg[15:8] == 132) || 
(freg[15:8] == 132 && treg[15:8] == 133) || 
(treg[15:8] == 132 && freg[15:8] == 133) || 
(freg[15:8] == 133 && treg[15:8] == 134) || 
(treg[15:8] == 133 && freg[15:8] == 134) || 
(freg[15:8] == 134 && treg[15:8] == 135) || 
(treg[15:8] == 134 && freg[15:8] == 135) || 
(freg[15:8] == 135 && treg[15:8] == 136) || 
(treg[15:8] == 135 && freg[15:8] == 136) || 
(freg[15:8] == 136 && treg[15:8] == 137) || 
(treg[15:8] == 136 && freg[15:8] == 137) || 
(freg[15:8] == 137 && treg[15:8] == 138) || 
(treg[15:8] == 137 && freg[15:8] == 138) || 
(freg[15:8] == 138 && treg[15:8] == 139) || 
(treg[15:8] == 138 && freg[15:8] == 139) || 
(freg[15:8] == 139 && treg[15:8] == 140) || 
(treg[15:8] == 139 && freg[15:8] == 140) || 
(freg[15:8] == 140 && treg[15:8] == 141) || 
(treg[15:8] == 140 && freg[15:8] == 141) || 
(freg[15:8] == 141 && treg[15:8] == 142) || 
(treg[15:8] == 141 && freg[15:8] == 142) || 
(freg[15:8] == 142 && treg[15:8] == 143) || 
(treg[15:8] == 142 && freg[15:8] == 143) || 
(freg[15:8] == 143 && treg[15:8] == 144) || 
(treg[15:8] == 143 && freg[15:8] == 144) || 
(freg[15:8] == 144 && treg[15:8] == 145) || 
(treg[15:8] == 144 && freg[15:8] == 145) || 
(freg[15:8] == 145 && treg[15:8] == 146) || 
(treg[15:8] == 145 && freg[15:8] == 146) || 
(freg[15:8] == 146 && treg[15:8] == 147) || 
(treg[15:8] == 146 && freg[15:8] == 147) || 
(freg[15:8] == 147 && treg[15:8] == 148) || 
(treg[15:8] == 147 && freg[15:8] == 148) || 
(freg[15:8] == 148 && treg[15:8] == 149) || 
(treg[15:8] == 148 && freg[15:8] == 149) || 
(freg[15:8] == 149 && treg[15:8] == 150) || 
(treg[15:8] == 149 && freg[15:8] == 150) || 
(freg[15:8] == 150 && treg[15:8] == 151) || 
(treg[15:8] == 150 && freg[15:8] == 151) || 
(freg[15:8] == 151 && treg[15:8] == 152) || 
(treg[15:8] == 151 && freg[15:8] == 152) || 
(freg[15:8] == 152 && treg[15:8] == 153) || 
(treg[15:8] == 152 && freg[15:8] == 153) || 
(freg[15:8] == 153 && treg[15:8] == 154) || 
(treg[15:8] == 153 && freg[15:8] == 154) || 
(freg[15:8] == 154 && treg[15:8] == 155) || 
(treg[15:8] == 154 && freg[15:8] == 155) || 
(freg[15:8] == 155 && treg[15:8] == 156) || 
(treg[15:8] == 155 && freg[15:8] == 156) || 
(freg[15:8] == 156 && treg[15:8] == 157) || 
(treg[15:8] == 156 && freg[15:8] == 157) || 
(freg[15:8] == 157 && treg[15:8] == 158) || 
(treg[15:8] == 157 && freg[15:8] == 158) || 
(freg[15:8] == 158 && treg[15:8] == 159) || 
(treg[15:8] == 158 && freg[15:8] == 159) || 
(freg[15:8] == 159 && treg[15:8] == 160) || 
(treg[15:8] == 159 && freg[15:8] == 160) || 
(freg[15:8] == 160 && treg[15:8] == 161) || 
(treg[15:8] == 160 && freg[15:8] == 161) || 
(freg[15:8] == 161 && treg[15:8] == 162) || 
(treg[15:8] == 161 && freg[15:8] == 162) || 
(freg[15:8] == 162 && treg[15:8] == 163) || 
(treg[15:8] == 162 && freg[15:8] == 163) || 
(freg[15:8] == 163 && treg[15:8] == 164) || 
(treg[15:8] == 163 && freg[15:8] == 164) || 
(freg[15:8] == 164 && treg[15:8] == 165) || 
(treg[15:8] == 164 && freg[15:8] == 165) || 
(freg[15:8] == 165 && treg[15:8] == 166) || 
(treg[15:8] == 165 && freg[15:8] == 166) || 
(freg[15:8] == 166 && treg[15:8] == 167) || 
(treg[15:8] == 166 && freg[15:8] == 167) || 
(freg[15:8] == 167 && treg[15:8] == 168) || 
(treg[15:8] == 167 && freg[15:8] == 168) || 
(freg[15:8] == 168 && treg[15:8] == 169) || 
(treg[15:8] == 168 && freg[15:8] == 169) || 
(freg[15:8] == 169 && treg[15:8] == 170) || 
(treg[15:8] == 169 && freg[15:8] == 170) || 
(freg[15:8] == 170 && treg[15:8] == 171) || 
(treg[15:8] == 170 && freg[15:8] == 171) || 
(freg[15:8] == 171 && treg[15:8] == 172) || 
(treg[15:8] == 171 && freg[15:8] == 172) || 
(freg[15:8] == 172 && treg[15:8] == 173) || 
(treg[15:8] == 172 && freg[15:8] == 173) || 
(freg[15:8] == 173 && treg[15:8] == 174) || 
(treg[15:8] == 173 && freg[15:8] == 174) || 
(freg[15:8] == 174 && treg[15:8] == 175) || 
(treg[15:8] == 174 && freg[15:8] == 175) || 
(freg[15:8] == 175 && treg[15:8] == 176) || 
(treg[15:8] == 175 && freg[15:8] == 176) || 
(freg[15:8] == 176 && treg[15:8] == 177) || 
(treg[15:8] == 176 && freg[15:8] == 177) || 
(freg[15:8] == 177 && treg[15:8] == 178) || 
(treg[15:8] == 177 && freg[15:8] == 178) || 
(freg[15:8] == 178 && treg[15:8] == 179) || 
(treg[15:8] == 178 && freg[15:8] == 179) || 
(freg[15:8] == 179 && treg[15:8] == 180) || 
(treg[15:8] == 179 && freg[15:8] == 180) || 
(freg[15:8] == 180 && treg[15:8] == 181) || 
(treg[15:8] == 180 && freg[15:8] == 181) || 
(freg[15:8] == 181 && treg[15:8] == 182) || 
(treg[15:8] == 181 && freg[15:8] == 182) || 
(freg[15:8] == 182 && treg[15:8] == 183) || 
(treg[15:8] == 182 && freg[15:8] == 183) || 
(freg[15:8] == 183 && treg[15:8] == 184) || 
(treg[15:8] == 183 && freg[15:8] == 184) || 
(freg[15:8] == 184 && treg[15:8] == 185) || 
(treg[15:8] == 184 && freg[15:8] == 185) || 
(freg[15:8] == 185 && treg[15:8] == 186) || 
(treg[15:8] == 185 && freg[15:8] == 186) || 
(freg[15:8] == 186 && treg[15:8] == 187) || 
(treg[15:8] == 186 && freg[15:8] == 187) || 
(freg[15:8] == 187 && treg[15:8] == 188) || 
(treg[15:8] == 187 && freg[15:8] == 188) || 
(freg[15:8] == 188 && treg[15:8] == 189) || 
(treg[15:8] == 188 && freg[15:8] == 189) || 
(freg[15:8] == 189 && treg[15:8] == 190) || 
(treg[15:8] == 189 && freg[15:8] == 190) || 
(freg[15:8] == 190 && treg[15:8] == 191) || 
(treg[15:8] == 190 && freg[15:8] == 191) || 
(freg[15:8] == 191 && treg[15:8] == 192) || 
(treg[15:8] == 191 && freg[15:8] == 192) || 
(freg[15:8] == 192 && treg[15:8] == 193) || 
(treg[15:8] == 192 && freg[15:8] == 193) || 
(freg[15:8] == 193 && treg[15:8] == 194) || 
(treg[15:8] == 193 && freg[15:8] == 194) || 
(freg[15:8] == 194 && treg[15:8] == 195) || 
(treg[15:8] == 194 && freg[15:8] == 195) || 
(freg[15:8] == 195 && treg[15:8] == 196) || 
(treg[15:8] == 195 && freg[15:8] == 196) || 
(freg[15:8] == 196 && treg[15:8] == 197) || 
(treg[15:8] == 196 && freg[15:8] == 197) || 
(freg[15:8] == 197 && treg[15:8] == 198) || 
(treg[15:8] == 197 && freg[15:8] == 198) || 
(freg[15:8] == 198 && treg[15:8] == 199) || 
(treg[15:8] == 198 && freg[15:8] == 199) || 
(freg[15:8] == 199 && treg[15:8] == 200) || 
(treg[15:8] == 199 && freg[15:8] == 200) || 
(freg[15:8] == 200 && treg[15:8] == 201) || 
(treg[15:8] == 200 && freg[15:8] == 201) || 
(freg[15:8] == 201 && treg[15:8] == 202) || 
(treg[15:8] == 201 && freg[15:8] == 202) || 
(freg[15:8] == 202 && treg[15:8] == 203) || 
(treg[15:8] == 202 && freg[15:8] == 203) || 
(freg[15:8] == 203 && treg[15:8] == 204) || 
(treg[15:8] == 203 && freg[15:8] == 204) || 
(freg[15:8] == 204 && treg[15:8] == 205) || 
(treg[15:8] == 204 && freg[15:8] == 205) || 
(freg[15:8] == 205 && treg[15:8] == 206) || 
(treg[15:8] == 205 && freg[15:8] == 206) || 
(freg[15:8] == 206 && treg[15:8] == 207) || 
(treg[15:8] == 206 && freg[15:8] == 207) || 
(freg[15:8] == 207 && treg[15:8] == 208) || 
(treg[15:8] == 207 && freg[15:8] == 208) || 
(freg[15:8] == 208 && treg[15:8] == 209) || 
(treg[15:8] == 208 && freg[15:8] == 209) || 
(freg[15:8] == 209 && treg[15:8] == 210) || 
(treg[15:8] == 209 && freg[15:8] == 210) || 
(freg[15:8] == 210 && treg[15:8] == 211) || 
(treg[15:8] == 210 && freg[15:8] == 211) || 
(freg[15:8] == 211 && treg[15:8] == 212) || 
(treg[15:8] == 211 && freg[15:8] == 212) || 
(freg[15:8] == 212 && treg[15:8] == 213) || 
(treg[15:8] == 212 && freg[15:8] == 213) || 
(freg[15:8] == 213 && treg[15:8] == 214) || 
(treg[15:8] == 213 && freg[15:8] == 214) || 
(freg[15:8] == 214 && treg[15:8] == 215) || 
(treg[15:8] == 214 && freg[15:8] == 215) || 
(freg[15:8] == 215 && treg[15:8] == 216) || 
(treg[15:8] == 215 && freg[15:8] == 216) || 
(freg[15:8] == 216 && treg[15:8] == 217) || 
(treg[15:8] == 216 && freg[15:8] == 217) || 
(freg[15:8] == 217 && treg[15:8] == 218) || 
(treg[15:8] == 217 && freg[15:8] == 218) || 
(freg[15:8] == 218 && treg[15:8] == 219) || 
(treg[15:8] == 218 && freg[15:8] == 219) || 
(freg[15:8] == 219 && treg[15:8] == 220) || 
(treg[15:8] == 219 && freg[15:8] == 220) || 
(freg[15:8] == 220 && treg[15:8] == 221) || 
(treg[15:8] == 220 && freg[15:8] == 221) || 
(freg[15:8] == 221 && treg[15:8] == 222) || 
(treg[15:8] == 221 && freg[15:8] == 222) || 
(freg[15:8] == 222 && treg[15:8] == 223) || 
(treg[15:8] == 222 && freg[15:8] == 223) || 
(freg[15:8] == 223 && treg[15:8] == 224) || 
(treg[15:8] == 223 && freg[15:8] == 224) || 
(freg[15:8] == 224 && treg[15:8] == 225) || 
(treg[15:8] == 224 && freg[15:8] == 225) || 
(freg[15:8] == 225 && treg[15:8] == 226) || 
(treg[15:8] == 225 && freg[15:8] == 226) || 
(freg[15:8] == 226 && treg[15:8] == 227) || 
(treg[15:8] == 226 && freg[15:8] == 227) || 
(freg[15:8] == 227 && treg[15:8] == 228) || 
(treg[15:8] == 227 && freg[15:8] == 228) || 
(freg[15:8] == 228 && treg[15:8] == 229) || 
(treg[15:8] == 228 && freg[15:8] == 229) || 
(freg[15:8] == 229 && treg[15:8] == 230) || 
(treg[15:8] == 229 && freg[15:8] == 230) || 
(freg[15:8] == 230 && treg[15:8] == 231) || 
(treg[15:8] == 230 && freg[15:8] == 231) || 
(freg[15:8] == 231 && treg[15:8] == 232) || 
(treg[15:8] == 231 && freg[15:8] == 232) || 
(freg[15:8] == 232 && treg[15:8] == 233) || 
(treg[15:8] == 232 && freg[15:8] == 233) || 
(freg[15:8] == 233 && treg[15:8] == 234) || 
(treg[15:8] == 233 && freg[15:8] == 234) || 
(freg[15:8] == 234 && treg[15:8] == 235) || 
(treg[15:8] == 234 && freg[15:8] == 235) || 
(freg[15:8] == 235 && treg[15:8] == 236) || 
(treg[15:8] == 235 && freg[15:8] == 236) || 
(freg[15:8] == 236 && treg[15:8] == 237) || 
(treg[15:8] == 236 && freg[15:8] == 237) || 
(freg[15:8] == 237 && treg[15:8] == 238) || 
(treg[15:8] == 237 && freg[15:8] == 238) || 
(freg[15:8] == 238 && treg[15:8] == 239) || 
(treg[15:8] == 238 && freg[15:8] == 239) || 
(freg[15:8] == 239 && treg[15:8] == 240) || 
(treg[15:8] == 239 && freg[15:8] == 240) || 
(freg[15:8] == 240 && treg[15:8] == 241) || 
(treg[15:8] == 240 && freg[15:8] == 241) || 
(freg[15:8] == 241 && treg[15:8] == 242) || 
(treg[15:8] == 241 && freg[15:8] == 242) || 
(freg[15:8] == 242 && treg[15:8] == 243) || 
(treg[15:8] == 242 && freg[15:8] == 243) || 
(freg[15:8] == 243 && treg[15:8] == 244) || 
(treg[15:8] == 243 && freg[15:8] == 244) || 
(freg[15:8] == 244 && treg[15:8] == 245) || 
(treg[15:8] == 244 && freg[15:8] == 245) || 
(freg[15:8] == 245 && treg[15:8] == 246) || 
(treg[15:8] == 245 && freg[15:8] == 246) || 
(freg[15:8] == 246 && treg[15:8] == 247) || 
(treg[15:8] == 246 && freg[15:8] == 247) || 
(freg[15:8] == 247 && treg[15:8] == 248) || 
(treg[15:8] == 247 && freg[15:8] == 248) || 
(freg[15:8] == 248 && treg[15:8] == 249) || 
(treg[15:8] == 248 && freg[15:8] == 249) || 
(freg[15:8] == 249 && treg[15:8] == 250) || 
(treg[15:8] == 249 && freg[15:8] == 250) || 
(freg[15:8] == 250 && treg[15:8] == 251) || 
(treg[15:8] == 250 && freg[15:8] == 251) || 
(freg[15:8] == 251 && treg[15:8] == 252) || 
(treg[15:8] == 251 && freg[15:8] == 252) || 
(freg[15:8] == 252 && treg[15:8] == 253) || 
(treg[15:8] == 252 && freg[15:8] == 253) || 
(freg[15:8] == 253 && treg[15:8] == 254) || 
(treg[15:8] == 253 && freg[15:8] == 254) || 
(freg[15:8] == 254 && treg[15:8] == 255) || 
(treg[15:8] == 254 && freg[15:8] == 255) || 
(freg[15:8] == 255 && treg[15:8] == 256) || 
(treg[15:8] == 255 && freg[15:8] == 256) || 
(freg[15:8] == 256 && treg[15:8] == 257) || 
(treg[15:8] == 256 && freg[15:8] == 257) || 
(freg[15:8] == 257 && treg[15:8] == 258) || 
(treg[15:8] == 257 && freg[15:8] == 258) || 
(freg[15:8] == 258 && treg[15:8] == 259) || 
(treg[15:8] == 258 && freg[15:8] == 259) || 
(freg[15:8] == 259 && treg[15:8] == 260) || 
(treg[15:8] == 259 && freg[15:8] == 260) || 
(freg[15:8] == 260 && treg[15:8] == 261) || 
(treg[15:8] == 260 && freg[15:8] == 261) || 
(freg[15:8] == 261 && treg[15:8] == 262) || 
(treg[15:8] == 261 && freg[15:8] == 262) || 
(freg[15:8] == 262 && treg[15:8] == 263) || 
(treg[15:8] == 262 && freg[15:8] == 263) || 
(freg[15:8] == 253 && treg[15:8] == 254) || 
(treg[15:8] == 253 && freg[15:8] == 254) || 
(freg[15:8] == 254 && treg[15:8] == 255) || 
(treg[15:8] == 254 && freg[15:8] == 255)
 
)                        
                    ||    //sliding within rows
                   (treg[11:6] == freg[11:6] && ((freg[7:0] == 0 && treg[7:0] == 1) || 
(treg[7:0] == 0 && freg[7:0] == 1) || 
(freg[7:0] == 1 && treg[7:0] == 2) || 
(treg[7:0] == 1 && freg[7:0] == 2) || 
(freg[7:0] == 2 && treg[7:0] == 3) || 
(treg[7:0] == 2 && freg[7:0] == 3) || 
(freg[7:0] == 3 && treg[7:0] == 4) || 
(treg[7:0] == 3 && freg[7:0] == 4) || 
(freg[7:0] == 4 && treg[7:0] == 5) || 
(treg[7:0] == 4 && freg[7:0] == 5) || 
(freg[7:0] == 5 && treg[7:0] == 6) || 
(treg[7:0] == 5 && freg[7:0] == 6) || 
(freg[7:0] == 6 && treg[7:0] == 7) || 
(treg[7:0] == 6 && freg[7:0] == 7) || 
(freg[7:0] == 7 && treg[7:0] == 8) || 
(treg[7:0] == 7 && freg[7:0] == 8) || 
(freg[7:0] == 8 && treg[7:0] == 9) || 
(treg[7:0] == 8 && freg[7:0] == 9) || 
(freg[7:0] == 9 && treg[7:0] == 10) || 
(treg[7:0] == 9 && freg[7:0] == 10) || 
(freg[7:0] == 10 && treg[7:0] == 11) || 
(treg[7:0] == 10 && freg[7:0] == 11) || 
(freg[7:0] == 11 && treg[7:0] == 12) || 
(treg[7:0] == 11 && freg[7:0] == 12) || 
(freg[7:0] == 12 && treg[7:0] == 13) || 
(treg[7:0] == 12 && freg[7:0] == 13) || 
(freg[7:0] == 13 && treg[7:0] == 14) || 
(treg[7:0] == 13 && freg[7:0] == 14) || 
(freg[7:0] == 14 && treg[7:0] == 15) || 
(treg[7:0] == 14 && freg[7:0] == 15) || 
(freg[7:0] == 15 && treg[7:0] == 16) || 
(treg[7:0] == 15 && freg[7:0] == 16) || 
(freg[7:0] == 16 && treg[7:0] == 17) || 
(treg[7:0] == 16 && freg[7:0] == 17) || 
(freg[7:0] == 17 && treg[7:0] == 18) || 
(treg[7:0] == 17 && freg[7:0] == 18) || 
(freg[7:0] == 18 && treg[7:0] == 19) || 
(treg[7:0] == 18 && freg[7:0] == 19) || 
(freg[7:0] == 19 && treg[7:0] == 20) || 
(treg[7:0] == 19 && freg[7:0] == 20) || 
(freg[7:0] == 20 && treg[7:0] == 21) || 
(treg[7:0] == 20 && freg[7:0] == 21) || 
(freg[7:0] == 21 && treg[7:0] == 22) || 
(treg[7:0] == 21 && freg[7:0] == 22) || 
(freg[7:0] == 22 && treg[7:0] == 23) || 
(treg[7:0] == 22 && freg[7:0] == 23) || 
(freg[7:0] == 23 && treg[7:0] == 24) || 
(treg[7:0] == 23 && freg[7:0] == 24) || 
(freg[7:0] == 24 && treg[7:0] == 25) || 
(treg[7:0] == 24 && freg[7:0] == 25) || 
(freg[7:0] == 25 && treg[7:0] == 26) || 
(treg[7:0] == 25 && freg[7:0] == 26) || 
(freg[7:0] == 26 && treg[7:0] == 27) || 
(treg[7:0] == 26 && freg[7:0] == 27) || 
(freg[7:0] == 27 && treg[7:0] == 28) || 
(treg[7:0] == 27 && freg[7:0] == 28) || 
(freg[7:0] == 28 && treg[7:0] == 29) || 
(treg[7:0] == 28 && freg[7:0] == 29) || 
(freg[7:0] == 29 && treg[7:0] == 30) || 
(treg[7:0] == 29 && freg[7:0] == 30) || 
(freg[7:0] == 30 && treg[7:0] == 31) || 
(treg[7:0] == 30 && freg[7:0] == 31) || 
(freg[7:0] == 31 && treg[7:0] == 32) || 
(treg[7:0] == 31 && freg[7:0] == 32) || 
(freg[7:0] == 32 && treg[7:0] == 33) || 
(treg[7:0] == 32 && freg[7:0] == 33) || 
(freg[7:0] == 33 && treg[7:0] == 34) || 
(treg[7:0] == 33 && freg[7:0] == 34) || 
(freg[7:0] == 34 && treg[7:0] == 35) || 
(treg[7:0] == 34 && freg[7:0] == 35) || 
(freg[7:0] == 35 && treg[7:0] == 36) || 
(treg[7:0] == 35 && freg[7:0] == 36) || 
(freg[7:0] == 36 && treg[7:0] == 37) || 
(treg[7:0] == 36 && freg[7:0] == 37) || 
(freg[7:0] == 37 && treg[7:0] == 38) || 
(treg[7:0] == 37 && freg[7:0] == 38) || 
(freg[7:0] == 38 && treg[7:0] == 39) || 
(treg[7:0] == 38 && freg[7:0] == 39) || 
(freg[7:0] == 39 && treg[7:0] == 40) || 
(treg[7:0] == 39 && freg[7:0] == 40) || 
(freg[7:0] == 40 && treg[7:0] == 41) || 
(treg[7:0] == 40 && freg[7:0] == 41) || 
(freg[7:0] == 41 && treg[7:0] == 42) || 
(treg[7:0] == 41 && freg[7:0] == 42) || 
(freg[7:0] == 42 && treg[7:0] == 43) || 
(treg[7:0] == 42 && freg[7:0] == 43) || 
(freg[7:0] == 43 && treg[7:0] == 44) || 
(treg[7:0] == 43 && freg[7:0] == 44) || 
(freg[7:0] == 44 && treg[7:0] == 45) || 
(treg[7:0] == 44 && freg[7:0] == 45) || 
(freg[7:0] == 45 && treg[7:0] == 46) || 
(treg[7:0] == 45 && freg[7:0] == 46) || 
(freg[7:0] == 46 && treg[7:0] == 47) || 
(treg[7:0] == 46 && freg[7:0] == 47) || 
(freg[7:0] == 47 && treg[7:0] == 48) || 
(treg[7:0] == 47 && freg[7:0] == 48) || 
(freg[7:0] == 48 && treg[7:0] == 49) || 
(treg[7:0] == 48 && freg[7:0] == 49) || 
(freg[7:0] == 49 && treg[7:0] == 50) || 
(treg[7:0] == 49 && freg[7:0] == 50) || 
(freg[7:0] == 50 && treg[7:0] == 51) || 
(treg[7:0] == 50 && freg[7:0] == 51) || 
(freg[7:0] == 51 && treg[7:0] == 52) || 
(treg[7:0] == 51 && freg[7:0] == 52) || 
(freg[7:0] == 52 && treg[7:0] == 53) || 
(treg[7:0] == 52 && freg[7:0] == 53) || 
(freg[7:0] == 53 && treg[7:0] == 54) || 
(treg[7:0] == 53 && freg[7:0] == 54) || 
(freg[7:0] == 54 && treg[7:0] == 55) || 
(treg[7:0] == 54 && freg[7:0] == 55) || 
(freg[7:0] == 55 && treg[7:0] == 56) || 
(treg[7:0] == 55 && freg[7:0] == 56) || 
(freg[7:0] == 56 && treg[7:0] == 57) || 
(treg[7:0] == 56 && freg[7:0] == 57) || 
(freg[7:0] == 57 && treg[7:0] == 58) || 
(treg[7:0] == 57 && freg[7:0] == 58) || 
(freg[7:0] == 58 && treg[7:0] == 59) || 
(treg[7:0] == 58 && freg[7:0] == 59) || 
(freg[7:0] == 59 && treg[7:0] == 60) || 
(treg[7:0] == 59 && freg[7:0] == 60) || 
(freg[7:0] == 60 && treg[7:0] == 61) || 
(treg[7:0] == 60 && freg[7:0] == 61) || 
(freg[7:0] == 61 && treg[7:0] == 62) || 
(treg[7:0] == 61 && freg[7:0] == 62) || 
(freg[7:0] == 62 && treg[7:0] == 63) || 
(treg[7:0] == 62 && freg[7:0] == 63) || 
(freg[7:0] == 63 && treg[7:0] == 64) || 
(treg[7:0] == 63 && freg[7:0] == 64) || 
(freg[7:0] == 64 && treg[7:0] == 65) || 
(treg[7:0] == 64 && freg[7:0] == 65) || 
(freg[7:0] == 65 && treg[7:0] == 66) || 
(treg[7:0] == 65 && freg[7:0] == 66) || 
(freg[7:0] == 66 && treg[7:0] == 67) || 
(treg[7:0] == 66 && freg[7:0] == 67) || 
(freg[7:0] == 67 && treg[7:0] == 68) || 
(treg[7:0] == 67 && freg[7:0] == 68) || 
(freg[7:0] == 68 && treg[7:0] == 69) || 
(treg[7:0] == 68 && freg[7:0] == 69) || 
(freg[7:0] == 69 && treg[7:0] == 70) || 
(treg[7:0] == 69 && freg[7:0] == 70) || 
(freg[7:0] == 70 && treg[7:0] == 71) || 
(treg[7:0] == 70 && freg[7:0] == 71) || 
(freg[7:0] == 71 && treg[7:0] == 72) || 
(treg[7:0] == 71 && freg[7:0] == 72) || 
(freg[7:0] == 72 && treg[7:0] == 73) || 
(treg[7:0] == 72 && freg[7:0] == 73) || 
(freg[7:0] == 73 && treg[7:0] == 74) || 
(treg[7:0] == 73 && freg[7:0] == 74) || 
(freg[7:0] == 74 && treg[7:0] == 75) || 
(treg[7:0] == 74 && freg[7:0] == 75) || 
(freg[7:0] == 75 && treg[7:0] == 76) || 
(treg[7:0] == 75 && freg[7:0] == 76) || 
(freg[7:0] == 76 && treg[7:0] == 77) || 
(treg[7:0] == 76 && freg[7:0] == 77) || 
(freg[7:0] == 77 && treg[7:0] == 78) || 
(treg[7:0] == 77 && freg[7:0] == 78) || 
(freg[7:0] == 78 && treg[7:0] == 79) || 
(treg[7:0] == 78 && freg[7:0] == 79) || 
(freg[7:0] == 79 && treg[7:0] == 80) || 
(treg[7:0] == 79 && freg[7:0] == 80) || 
(freg[7:0] == 80 && treg[7:0] == 81) || 
(treg[7:0] == 80 && freg[7:0] == 81) || 
(freg[7:0] == 81 && treg[7:0] == 82) || 
(treg[7:0] == 81 && freg[7:0] == 82) || 
(freg[7:0] == 82 && treg[7:0] == 83) || 
(treg[7:0] == 82 && freg[7:0] == 83) || 
(freg[7:0] == 83 && treg[7:0] == 84) || 
(treg[7:0] == 83 && freg[7:0] == 84) || 
(freg[7:0] == 84 && treg[7:0] == 85) || 
(treg[7:0] == 84 && freg[7:0] == 85) || 
(freg[7:0] == 85 && treg[7:0] == 86) || 
(treg[7:0] == 85 && freg[7:0] == 86) || 
(freg[7:0] == 86 && treg[7:0] == 87) || 
(treg[7:0] == 86 && freg[7:0] == 87) || 
(freg[7:0] == 87 && treg[7:0] == 88) || 
(treg[7:0] == 87 && freg[7:0] == 88) || 
(freg[7:0] == 88 && treg[7:0] == 89) || 
(treg[7:0] == 88 && freg[7:0] == 89) || 
(freg[7:0] == 89 && treg[7:0] == 90) || 
(treg[7:0] == 89 && freg[7:0] == 90) || 
(freg[7:0] == 90 && treg[7:0] == 91) || 
(treg[7:0] == 90 && freg[7:0] == 91) || 
(freg[7:0] == 91 && treg[7:0] == 92) || 
(treg[7:0] == 91 && freg[7:0] == 92) || 
(freg[7:0] == 92 && treg[7:0] == 93) || 
(treg[7:0] == 92 && freg[7:0] == 93) || 
(freg[7:0] == 93 && treg[7:0] == 94) || 
(treg[7:0] == 93 && freg[7:0] == 94) || 
(freg[7:0] == 94 && treg[7:0] == 95) || 
(treg[7:0] == 94 && freg[7:0] == 95) || 
(freg[7:0] == 95 && treg[7:0] == 96) || 
(treg[7:0] == 95 && freg[7:0] == 96) || 
(freg[7:0] == 96 && treg[7:0] == 97) || 
(treg[7:0] == 96 && freg[7:0] == 97) || 
(freg[7:0] == 97 && treg[7:0] == 98) || 
(treg[7:0] == 97 && freg[7:0] == 98) || 
(freg[7:0] == 98 && treg[7:0] == 99) || 
(treg[7:0] == 98 && freg[7:0] == 99) || 
(freg[7:0] == 99 && treg[7:0] == 100) || 
(treg[7:0] == 99 && freg[7:0] == 100) || 
(freg[7:0] == 100 && treg[7:0] == 101) || 
(treg[7:0] == 100 && freg[7:0] == 101) || 
(freg[7:0] == 101 && treg[7:0] == 102) || 
(treg[7:0] == 101 && freg[7:0] == 102) || 
(freg[7:0] == 102 && treg[7:0] == 103) || 
(treg[7:0] == 102 && freg[7:0] == 103) || 
(freg[7:0] == 103 && treg[7:0] == 104) || 
(treg[7:0] == 103 && freg[7:0] == 104) || 
(freg[7:0] == 104 && treg[7:0] == 105) || 
(treg[7:0] == 104 && freg[7:0] == 105) || 
(freg[7:0] == 105 && treg[7:0] == 106) || 
(treg[7:0] == 105 && freg[7:0] == 106) || 
(freg[7:0] == 106 && treg[7:0] == 107) || 
(treg[7:0] == 106 && freg[7:0] == 107) || 
(freg[7:0] == 107 && treg[7:0] == 108) || 
(treg[7:0] == 107 && freg[7:0] == 108) || 
(freg[7:0] == 108 && treg[7:0] == 109) || 
(treg[7:0] == 108 && freg[7:0] == 109) || 
(freg[7:0] == 109 && treg[7:0] == 110) || 
(treg[7:0] == 109 && freg[7:0] == 110) || 
(freg[7:0] == 110 && treg[7:0] == 111) || 
(treg[7:0] == 110 && freg[7:0] == 111) || 
(freg[7:0] == 111 && treg[7:0] == 112) || 
(treg[7:0] == 111 && freg[7:0] == 112) || 
(freg[7:0] == 112 && treg[7:0] == 113) || 
(treg[7:0] == 112 && freg[7:0] == 113) || 
(freg[7:0] == 113 && treg[7:0] == 114) || 
(treg[7:0] == 113 && freg[7:0] == 114) || 
(freg[7:0] == 114 && treg[7:0] == 115) || 
(treg[7:0] == 114 && freg[7:0] == 115) || 
(freg[7:0] == 115 && treg[7:0] == 116) || 
(treg[7:0] == 115 && freg[7:0] == 116) || 
(freg[7:0] == 116 && treg[7:0] == 117) || 
(treg[7:0] == 116 && freg[7:0] == 117) || 
(freg[7:0] == 117 && treg[7:0] == 118) || 
(treg[7:0] == 117 && freg[7:0] == 118) || 
(freg[7:0] == 118 && treg[7:0] == 119) || 
(treg[7:0] == 118 && freg[7:0] == 119) || 
(freg[7:0] == 119 && treg[7:0] == 120) || 
(treg[7:0] == 119 && freg[7:0] == 120) || 
(freg[7:0] == 120 && treg[7:0] == 121) || 
(treg[7:0] == 120 && freg[7:0] == 121) || 
(freg[7:0] == 121 && treg[7:0] == 122) || 
(treg[7:0] == 121 && freg[7:0] == 122) || 
(freg[7:0] == 122 && treg[7:0] == 123) || 
(treg[7:0] == 122 && freg[7:0] == 123) || 
(freg[7:0] == 123 && treg[7:0] == 124) || 
(treg[7:0] == 123 && freg[7:0] == 124) || 
(freg[7:0] == 124 && treg[7:0] == 125) || 
(treg[7:0] == 124 && freg[7:0] == 125) || 
(freg[7:0] == 125 && treg[7:0] == 126) || 
(treg[7:0] == 125 && freg[7:0] == 126) || 
(freg[7:0] == 126 && treg[7:0] == 127) || 
(treg[7:0] == 126 && freg[7:0] == 127) || 
(freg[7:0] == 127 && treg[7:0] == 128) || 
(treg[7:0] == 127 && freg[7:0] == 128) || 
(freg[7:0] == 128 && treg[7:0] == 129) || 
(treg[7:0] == 128 && freg[7:0] == 129) || 
(freg[7:0] == 129 && treg[7:0] == 130) || 
(treg[7:0] == 129 && freg[7:0] == 130) || 
(freg[7:0] == 130 && treg[7:0] == 131) || 
(treg[7:0] == 130 && freg[7:0] == 131) || 
(freg[7:0] == 131 && treg[7:0] == 132) || 
(treg[7:0] == 131 && freg[7:0] == 132) || 
(freg[7:0] == 132 && treg[7:0] == 133) || 
(treg[7:0] == 132 && freg[7:0] == 133) || 
(freg[7:0] == 133 && treg[7:0] == 134) || 
(treg[7:0] == 133 && freg[7:0] == 134) || 
(freg[7:0] == 134 && treg[7:0] == 135) || 
(treg[7:0] == 134 && freg[7:0] == 135) || 
(freg[7:0] == 135 && treg[7:0] == 136) || 
(treg[7:0] == 135 && freg[7:0] == 136) || 
(freg[7:0] == 136 && treg[7:0] == 137) || 
(treg[7:0] == 136 && freg[7:0] == 137) || 
(freg[7:0] == 137 && treg[7:0] == 138) || 
(treg[7:0] == 137 && freg[7:0] == 138) || 
(freg[7:0] == 138 && treg[7:0] == 139) || 
(treg[7:0] == 138 && freg[7:0] == 139) || 
(freg[7:0] == 139 && treg[7:0] == 140) || 
(treg[7:0] == 139 && freg[7:0] == 140) || 
(freg[7:0] == 140 && treg[7:0] == 141) || 
(treg[7:0] == 140 && freg[7:0] == 141) || 
(freg[7:0] == 141 && treg[7:0] == 142) || 
(treg[7:0] == 141 && freg[7:0] == 142) || 
(freg[7:0] == 142 && treg[7:0] == 143) || 
(treg[7:0] == 142 && freg[7:0] == 143) || 
(freg[7:0] == 143 && treg[7:0] == 144) || 
(treg[7:0] == 143 && freg[7:0] == 144) || 
(freg[7:0] == 144 && treg[7:0] == 145) || 
(treg[7:0] == 144 && freg[7:0] == 145) || 
(freg[7:0] == 145 && treg[7:0] == 146) || 
(treg[7:0] == 145 && freg[7:0] == 146) || 
(freg[7:0] == 146 && treg[7:0] == 147) || 
(treg[7:0] == 146 && freg[7:0] == 147) || 
(freg[7:0] == 147 && treg[7:0] == 148) || 
(treg[7:0] == 147 && freg[7:0] == 148) || 
(freg[7:0] == 148 && treg[7:0] == 149) || 
(treg[7:0] == 148 && freg[7:0] == 149) || 
(freg[7:0] == 149 && treg[7:0] == 150) || 
(treg[7:0] == 149 && freg[7:0] == 150) || 
(freg[7:0] == 150 && treg[7:0] == 151) || 
(treg[7:0] == 150 && freg[7:0] == 151) || 
(freg[7:0] == 151 && treg[7:0] == 152) || 
(treg[7:0] == 151 && freg[7:0] == 152) || 
(freg[7:0] == 152 && treg[7:0] == 153) || 
(treg[7:0] == 152 && freg[7:0] == 153) || 
(freg[7:0] == 153 && treg[7:0] == 154) || 
(treg[7:0] == 153 && freg[7:0] == 154) || 
(freg[7:0] == 154 && treg[7:0] == 155) || 
(treg[7:0] == 154 && freg[7:0] == 155) || 
(freg[7:0] == 155 && treg[7:0] == 156) || 
(treg[7:0] == 155 && freg[7:0] == 156) || 
(freg[7:0] == 156 && treg[7:0] == 157) || 
(treg[7:0] == 156 && freg[7:0] == 157) || 
(freg[7:0] == 157 && treg[7:0] == 158) || 
(treg[7:0] == 157 && freg[7:0] == 158) || 
(freg[7:0] == 158 && treg[7:0] == 159) || 
(treg[7:0] == 158 && freg[7:0] == 159) || 
(freg[7:0] == 159 && treg[7:0] == 160) || 
(treg[7:0] == 159 && freg[7:0] == 160) || 
(freg[7:0] == 160 && treg[7:0] == 161) || 
(treg[7:0] == 160 && freg[7:0] == 161) || 
(freg[7:0] == 161 && treg[7:0] == 162) || 
(treg[7:0] == 161 && freg[7:0] == 162) || 
(freg[7:0] == 162 && treg[7:0] == 163) || 
(treg[7:0] == 162 && freg[7:0] == 163) || 
(freg[7:0] == 163 && treg[7:0] == 164) || 
(treg[7:0] == 163 && freg[7:0] == 164) || 
(freg[7:0] == 164 && treg[7:0] == 165) || 
(treg[7:0] == 164 && freg[7:0] == 165) || 
(freg[7:0] == 165 && treg[7:0] == 166) || 
(treg[7:0] == 165 && freg[7:0] == 166) || 
(freg[7:0] == 166 && treg[7:0] == 167) || 
(treg[7:0] == 166 && freg[7:0] == 167) || 
(freg[7:0] == 167 && treg[7:0] == 168) || 
(treg[7:0] == 167 && freg[7:0] == 168) || 
(freg[7:0] == 168 && treg[7:0] == 169) || 
(treg[7:0] == 168 && freg[7:0] == 169) || 
(freg[7:0] == 169 && treg[7:0] == 170) || 
(treg[7:0] == 169 && freg[7:0] == 170) || 
(freg[7:0] == 170 && treg[7:0] == 171) || 
(treg[7:0] == 170 && freg[7:0] == 171) || 
(freg[7:0] == 171 && treg[7:0] == 172) || 
(treg[7:0] == 171 && freg[7:0] == 172) || 
(freg[7:0] == 172 && treg[7:0] == 173) || 
(treg[7:0] == 172 && freg[7:0] == 173) || 
(freg[7:0] == 173 && treg[7:0] == 174) || 
(treg[7:0] == 173 && freg[7:0] == 174) || 
(freg[7:0] == 174 && treg[7:0] == 175) || 
(treg[7:0] == 174 && freg[7:0] == 175) || 
(freg[7:0] == 175 && treg[7:0] == 176) || 
(treg[7:0] == 175 && freg[7:0] == 176) || 
(freg[7:0] == 176 && treg[7:0] == 177) || 
(treg[7:0] == 176 && freg[7:0] == 177) || 
(freg[7:0] == 177 && treg[7:0] == 178) || 
(treg[7:0] == 177 && freg[7:0] == 178) || 
(freg[7:0] == 178 && treg[7:0] == 179) || 
(treg[7:0] == 178 && freg[7:0] == 179) || 
(freg[7:0] == 179 && treg[7:0] == 180) || 
(treg[7:0] == 179 && freg[7:0] == 180) || 
(freg[7:0] == 180 && treg[7:0] == 181) || 
(treg[7:0] == 180 && freg[7:0] == 181) || 
(freg[7:0] == 181 && treg[7:0] == 182) || 
(treg[7:0] == 181 && freg[7:0] == 182) || 
(freg[7:0] == 182 && treg[7:0] == 183) || 
(treg[7:0] == 182 && freg[7:0] == 183) || 
(freg[7:0] == 183 && treg[7:0] == 184) || 
(treg[7:0] == 183 && freg[7:0] == 184) || 
(freg[7:0] == 184 && treg[7:0] == 185) || 
(treg[7:0] == 184 && freg[7:0] == 185) || 
(freg[7:0] == 185 && treg[7:0] == 186) || 
(treg[7:0] == 185 && freg[7:0] == 186) || 
(freg[7:0] == 186 && treg[7:0] == 187) || 
(treg[7:0] == 186 && freg[7:0] == 187) || 
(freg[7:0] == 187 && treg[7:0] == 188) || 
(treg[7:0] == 187 && freg[7:0] == 188) || 
(freg[7:0] == 188 && treg[7:0] == 189) || 
(treg[7:0] == 188 && freg[7:0] == 189) || 
(freg[7:0] == 189 && treg[7:0] == 190) || 
(treg[7:0] == 189 && freg[7:0] == 190) || 
(freg[7:0] == 190 && treg[7:0] == 191) || 
(treg[7:0] == 190 && freg[7:0] == 191) || 
(freg[7:0] == 191 && treg[7:0] == 192) || 
(treg[7:0] == 191 && freg[7:0] == 192) || 
(freg[7:0] == 192 && treg[7:0] == 193) || 
(treg[7:0] == 192 && freg[7:0] == 193) || 
(freg[7:0] == 193 && treg[7:0] == 194) || 
(treg[7:0] == 193 && freg[7:0] == 194) || 
(freg[7:0] == 194 && treg[7:0] == 195) || 
(treg[7:0] == 194 && freg[7:0] == 195) || 
(freg[7:0] == 195 && treg[7:0] == 196) || 
(treg[7:0] == 195 && freg[7:0] == 196) || 
(freg[7:0] == 196 && treg[7:0] == 197) || 
(treg[7:0] == 196 && freg[7:0] == 197) || 
(freg[7:0] == 197 && treg[7:0] == 198) || 
(treg[7:0] == 197 && freg[7:0] == 198) || 
(freg[7:0] == 198 && treg[7:0] == 199) || 
(treg[7:0] == 198 && freg[7:0] == 199) || 
(freg[7:0] == 199 && treg[7:0] == 200) || 
(treg[7:0] == 199 && freg[7:0] == 200) || 
(freg[7:0] == 200 && treg[7:0] == 201) || 
(treg[7:0] == 200 && freg[7:0] == 201) || 
(freg[7:0] == 201 && treg[7:0] == 202) || 
(treg[7:0] == 201 && freg[7:0] == 202) || 
(freg[7:0] == 202 && treg[7:0] == 203) || 
(treg[7:0] == 202 && freg[7:0] == 203) || 
(freg[7:0] == 203 && treg[7:0] == 204) || 
(treg[7:0] == 203 && freg[7:0] == 204) || 
(freg[7:0] == 204 && treg[7:0] == 205) || 
(treg[7:0] == 204 && freg[7:0] == 205) || 
(freg[7:0] == 205 && treg[7:0] == 206) || 
(treg[7:0] == 205 && freg[7:0] == 206) || 
(freg[7:0] == 206 && treg[7:0] == 207) || 
(treg[7:0] == 206 && freg[7:0] == 207) || 
(freg[7:0] == 207 && treg[7:0] == 208) || 
(treg[7:0] == 207 && freg[7:0] == 208) || 
(freg[7:0] == 208 && treg[7:0] == 209) || 
(treg[7:0] == 208 && freg[7:0] == 209) || 
(freg[7:0] == 209 && treg[7:0] == 210) || 
(treg[7:0] == 209 && freg[7:0] == 210) || 
(freg[7:0] == 210 && treg[7:0] == 211) || 
(treg[7:0] == 210 && freg[7:0] == 211) || 
(freg[7:0] == 211 && treg[7:0] == 212) || 
(treg[7:0] == 211 && freg[7:0] == 212) || 
(freg[7:0] == 212 && treg[7:0] == 213) || 
(treg[7:0] == 212 && freg[7:0] == 213) || 
(freg[7:0] == 213 && treg[7:0] == 214) || 
(treg[7:0] == 213 && freg[7:0] == 214) || 
(freg[7:0] == 214 && treg[7:0] == 215) || 
(treg[7:0] == 214 && freg[7:0] == 215) || 
(freg[7:0] == 215 && treg[7:0] == 216) || 
(treg[7:0] == 215 && freg[7:0] == 216) || 
(freg[7:0] == 216 && treg[7:0] == 217) || 
(treg[7:0] == 216 && freg[7:0] == 217) || 
(freg[7:0] == 217 && treg[7:0] == 218) || 
(treg[7:0] == 217 && freg[7:0] == 218) || 
(freg[7:0] == 218 && treg[7:0] == 219) || 
(treg[7:0] == 218 && freg[7:0] == 219) || 
(freg[7:0] == 219 && treg[7:0] == 220) || 
(treg[7:0] == 219 && freg[7:0] == 220) || 
(freg[7:0] == 220 && treg[7:0] == 221) || 
(treg[7:0] == 220 && freg[7:0] == 221) || 
(freg[7:0] == 221 && treg[7:0] == 222) || 
(treg[7:0] == 221 && freg[7:0] == 222) || 
(freg[7:0] == 222 && treg[7:0] == 223) || 
(treg[7:0] == 222 && freg[7:0] == 223) || 
(freg[7:0] == 223 && treg[7:0] == 224) || 
(treg[7:0] == 223 && freg[7:0] == 224) || 
(freg[7:0] == 224 && treg[7:0] == 225) || 
(treg[7:0] == 224 && freg[7:0] == 225) || 
(freg[7:0] == 225 && treg[7:0] == 226) || 
(treg[7:0] == 225 && freg[7:0] == 226) || 
(freg[7:0] == 226 && treg[7:0] == 227) || 
(treg[7:0] == 226 && freg[7:0] == 227) || 
(freg[7:0] == 227 && treg[7:0] == 228) || 
(treg[7:0] == 227 && freg[7:0] == 228) || 
(freg[7:0] == 228 && treg[7:0] == 229) || 
(treg[7:0] == 228 && freg[7:0] == 229) || 
(freg[7:0] == 229 && treg[7:0] == 230) || 
(treg[7:0] == 229 && freg[7:0] == 230) || 
(freg[7:0] == 230 && treg[7:0] == 231) || 
(treg[7:0] == 230 && freg[7:0] == 231) || 
(freg[7:0] == 231 && treg[7:0] == 232) || 
(treg[7:0] == 231 && freg[7:0] == 232) || 
(freg[7:0] == 232 && treg[7:0] == 233) || 
(treg[7:0] == 232 && freg[7:0] == 233) || 
(freg[7:0] == 233 && treg[7:0] == 234) || 
(treg[7:0] == 233 && freg[7:0] == 234) || 
(freg[7:0] == 234 && treg[7:0] == 235) || 
(treg[7:0] == 234 && freg[7:0] == 235) || 
(freg[7:0] == 235 && treg[7:0] == 236) || 
(treg[7:0] == 235 && freg[7:0] == 236) || 
(freg[7:0] == 236 && treg[7:0] == 237) || 
(treg[7:0] == 236 && freg[7:0] == 237) || 
(freg[7:0] == 237 && treg[7:0] == 238) || 
(treg[7:0] == 237 && freg[7:0] == 238) || 
(freg[7:0] == 238 && treg[7:0] == 239) || 
(treg[7:0] == 238 && freg[7:0] == 239) || 
(freg[7:0] == 239 && treg[7:0] == 240) || 
(treg[7:0] == 239 && freg[7:0] == 240) || 
(freg[7:0] == 240 && treg[7:0] == 241) || 
(treg[7:0] == 240 && freg[7:0] == 241) || 
(freg[7:0] == 241 && treg[7:0] == 242) || 
(treg[7:0] == 241 && freg[7:0] == 242) || 
(freg[7:0] == 242 && treg[7:0] == 243) || 
(treg[7:0] == 242 && freg[7:0] == 243) || 
(freg[7:0] == 243 && treg[7:0] == 244) || 
(treg[7:0] == 243 && freg[7:0] == 244) || 
(freg[7:0] == 244 && treg[7:0] == 245) || 
(treg[7:0] == 244 && freg[7:0] == 245) || 
(freg[7:0] == 245 && treg[7:0] == 246) || 
(treg[7:0] == 245 && freg[7:0] == 246) || 
(freg[7:0] == 246 && treg[7:0] == 247) || 
(treg[7:0] == 246 && freg[7:0] == 247) || 
(freg[7:0] == 247 && treg[7:0] == 248) || 
(treg[7:0] == 247 && freg[7:0] == 248) || 
(freg[7:0] == 248 && treg[7:0] == 249) || 
(treg[7:0] == 248 && freg[7:0] == 249) || 
(freg[7:0] == 249 && treg[7:0] == 250) || 
(treg[7:0] == 249 && freg[7:0] == 250) || 
(freg[7:0] == 250 && treg[7:0] == 251) || 
(treg[7:0] == 250 && freg[7:0] == 251) || 
(freg[7:0] == 251 && treg[7:0] == 252) || 
(treg[7:0] == 251 && freg[7:0] == 252) || 
(freg[7:0] == 252 && treg[7:0] == 253) || 
(treg[7:0] == 252 && freg[7:0] == 253) || 
(freg[7:0] == 253 && treg[7:0] == 254) || 
(treg[7:0] == 253 && freg[7:0] == 254) || 
(freg[7:0] == 254 && treg[7:0] == 255) || 
(treg[7:0] == 254 && freg[7:0] == 255)

 )))
                     );
    assign parity = 
	   (((b[0] & 5) == 1) | ((b[0] & 5) == 4)) ^
	   (((b[1] & 5) == 0) | ((b[1] & 5) == 5)) ^
	   (((b[2] & 5) == 1) | ((b[2] & 5) == 4)) ^
	   (((b[3] & 5) == 0) | ((b[3] & 5) == 5)) ^
	   (((b[4] & 5) == 1) | ((b[4] & 5) == 4)) ^
	   (((b[5] & 5) == 0) | ((b[5] & 5) == 5)) ^
	   (((b[6] & 5) == 1) | ((b[6] & 5) == 4)) ^
	   (((b[7] & 5) == 0) | ((b[7] & 5) == 5));
 
    always @(posedge clock) begin
	freg <= from;
	treg <= to;
    end

    always @(posedge clock) begin
	if (valid) begin
	    b[treg] <= b[freg];
	    b[freg] <= 0;
	end
    end

/*invariant property
!(b<*0*>[2:0]=0 * b<*1*>[2:0]=1 * b<*2*>[2:0]=2 * b<*3*>[2:0]=3 *
  b<*4*>[2:0]=4 * b<*5*>[2:0]=5 * b<*6*>[2:0]=6 * b<*7*>[2:0]=7);*/
	assert property (!(b[0] == 0 && 
b[1] == 1 && 
b[2] == 2 && 
b[3] == 3 && 
b[4] == 4 && 
b[5] == 5 && 
b[6] == 6 && 
b[7] == 7 && 
b[8] == 8 && 
b[9] == 9 && 
b[10] == 10 && 
b[11] == 11 && 
b[12] == 12 && 
b[13] == 13 && 
b[14] == 14 && 
b[15] == 15 && 
b[16] == 16 && 
b[17] == 17 && 
b[18] == 18 && 
b[19] == 19 && 
b[20] == 20 && 
b[21] == 21 && 
b[22] == 22 && 
b[23] == 23 && 
b[24] == 24 && 
b[25] == 25 && 
b[26] == 26 && 
b[27] == 27 && 
b[28] == 28 && 
b[29] == 29 && 
b[30] == 30 && 
b[31] == 31 && 
b[32] == 32 && 
b[33] == 33 && 
b[34] == 34 && 
b[35] == 35 && 
b[36] == 36 && 
b[37] == 37 && 
b[38] == 38 && 
b[39] == 39 && 
b[40] == 40 && 
b[41] == 41 && 
b[42] == 42 && 
b[43] == 43 && 
b[44] == 44 && 
b[45] == 45 && 
b[46] == 46 && 
b[47] == 47 && 
b[48] == 48 && 
b[49] == 49 && 
b[50] == 50 && 
b[51] == 51 && 
b[52] == 52 && 
b[53] == 53 && 
b[54] == 54 && 
b[55] == 55 && 
b[56] == 56 && 
b[57] == 57 && 
b[58] == 58 && 
b[59] == 59 && 
b[60] == 60 && 
b[61] == 61 && 
b[62] == 62 && 
b[63] == 63 && 
b[64] == 64 && 
b[65] == 65 && 
b[66] == 66 && 
b[67] == 67 && 
b[68] == 68 && 
b[69] == 69 && 
b[70] == 70 && 
b[71] == 71 && 
b[72] == 72 && 
b[73] == 73 && 
b[74] == 74 && 
b[75] == 75 && 
b[76] == 76 && 
b[77] == 77 && 
b[78] == 78 && 
b[79] == 79 && 
b[80] == 80 && 
b[81] == 81 && 
b[82] == 82 && 
b[83] == 83 && 
b[84] == 84 && 
b[85] == 85 && 
b[86] == 86 && 
b[87] == 87 && 
b[88] == 88 && 
b[89] == 89 && 
b[90] == 90 && 
b[91] == 91 && 
b[92] == 92 && 
b[93] == 93 && 
b[94] == 94 && 
b[95] == 95 && 
b[96] == 96 && 
b[97] == 97 && 
b[98] == 98 && 
b[99] == 99 && 
b[100] == 100 && 
b[101] == 101 && 
b[102] == 102 && 
b[103] == 103 && 
b[104] == 104 && 
b[105] == 105 && 
b[106] == 106 && 
b[107] == 107 && 
b[108] == 108 && 
b[109] == 109 && 
b[110] == 110 && 
b[111] == 111 && 
b[112] == 112 && 
b[113] == 113 && 
b[114] == 114 && 
b[115] == 115 && 
b[116] == 116 && 
b[117] == 117 && 
b[118] == 118 && 
b[119] == 119 && 
b[120] == 120 && 
b[121] == 121 && 
b[122] == 122 && 
b[123] == 123 && 
b[124] == 124 && 
b[125] == 125 && 
b[126] == 126 && 
b[127] == 127 && 
b[128] == 128 && 
b[129] == 129 && 
b[130] == 130 && 
b[131] == 131 && 
b[132] == 132 && 
b[133] == 133 && 
b[134] == 134 && 
b[135] == 135 && 
b[136] == 136 && 
b[137] == 137 && 
b[138] == 138 && 
b[139] == 139 && 
b[140] == 140 && 
b[141] == 141 && 
b[142] == 142 && 
b[143] == 143 && 
b[144] == 144 && 
b[145] == 145 && 
b[146] == 146 && 
b[147] == 147 && 
b[148] == 148 && 
b[149] == 149 && 
b[150] == 150 && 
b[151] == 151 && 
b[152] == 152 && 
b[153] == 153 && 
b[154] == 154 && 
b[155] == 155 && 
b[156] == 156 && 
b[157] == 157 && 
b[158] == 158 && 
b[159] == 159 && 
b[160] == 160 && 
b[161] == 161 && 
b[162] == 162 && 
b[163] == 163 && 
b[164] == 164 && 
b[165] == 165 && 
b[166] == 166 && 
b[167] == 167 && 
b[168] == 168 && 
b[169] == 169 && 
b[170] == 170 && 
b[171] == 171 && 
b[172] == 172 && 
b[173] == 173 && 
b[174] == 174 && 
b[175] == 175 && 
b[176] == 176 && 
b[177] == 177 && 
b[178] == 178 && 
b[179] == 179 && 
b[180] == 180 && 
b[181] == 181 && 
b[182] == 182 && 
b[183] == 183 && 
b[184] == 184 && 
b[185] == 185 && 
b[186] == 186 && 
b[187] == 187 && 
b[188] == 188 && 
b[189] == 189 && 
b[190] == 190 && 
b[191] == 191 && 
b[192] == 192 && 
b[193] == 193 && 
b[194] == 194 && 
b[195] == 195 && 
b[196] == 196 && 
b[197] == 197 && 
b[198] == 198 && 
b[199] == 199 && 
b[200] == 200 && 
b[201] == 201 && 
b[202] == 202 && 
b[203] == 203 && 
b[204] == 204 && 
b[205] == 205 && 
b[206] == 206 && 
b[207] == 207 && 
b[208] == 208 && 
b[209] == 209 && 
b[210] == 210 && 
b[211] == 211 && 
b[212] == 212 && 
b[213] == 213 && 
b[214] == 214 && 
b[215] == 215 && 
b[216] == 216 && 
b[217] == 217 && 
b[218] == 218 && 
b[219] == 219 && 
b[220] == 220 && 
b[221] == 221 && 
b[222] == 222 && 
b[223] == 223 && 
b[224] == 224 && 
b[225] == 225 && 
b[226] == 226 && 
b[227] == 227 && 
b[228] == 228 && 
b[229] == 229 && 
b[230] == 230 && 
b[231] == 231 && 
b[232] == 232 && 
b[233] == 233 && 
b[234] == 234 && 
b[235] == 235 && 
b[236] == 236 && 
b[237] == 237 && 
b[238] == 238 && 
b[239] == 239 && 
b[240] == 240 && 
b[241] == 241 && 
b[242] == 242 && 
b[243] == 243 && 
b[244] == 244 && 
b[245] == 245 && 
b[246] == 246 && 
b[247] == 247 && 
b[248] == 248 && 
b[249] == 249 && 
b[250] == 250 && 
b[251] == 251 && 
b[252] == 252 && 
b[253] == 253 && 
b[254] == 254 && 
b[255] == 255 && 
b[256] == 256 && 
b[257] == 257 && 
b[258] == 258 && 
b[259] == 259 && 
b[260] == 260 && 
b[261] == 261 && 
b[262] == 262 && 
b[263] == 263 && 
b[264] == 264 && 
b[265] == 265 && 
b[266] == 266 && 
b[267] == 267 && 
b[268] == 268 && 
b[269] == 269 && 
b[270] == 270 && 
b[271] == 271 && 
b[272] == 272 && 
b[273] == 273 && 
b[274] == 274 && 
b[275] == 275 && 
b[276] == 276 && 
b[277] == 277 && 
b[278] == 278 && 
b[279] == 279 && 
b[280] == 280 && 
b[281] == 281 && 
b[282] == 282 && 
b[283] == 283 && 
b[284] == 284 && 
b[285] == 285 && 
b[286] == 286 && 
b[287] == 287 && 
b[288] == 288 && 
b[289] == 289 && 
b[290] == 290 && 
b[291] == 291 && 
b[292] == 292 && 
b[293] == 293 && 
b[294] == 294 && 
b[295] == 295 && 
b[296] == 296 && 
b[297] == 297 && 
b[298] == 298 && 
b[299] == 299 && 
b[300] == 300 && 
b[301] == 301 && 
b[302] == 302 && 
b[303] == 303 && 
b[304] == 304 && 
b[305] == 305 && 
b[306] == 306 && 
b[307] == 307 && 
b[308] == 308 && 
b[309] == 309 && 
b[310] == 310 && 
b[311] == 311 && 
b[312] == 312 && 
b[313] == 313 && 
b[314] == 314 && 
b[315] == 315 && 
b[316] == 316 && 
b[317] == 317 && 
b[318] == 318 && 
b[319] == 319 && 
b[320] == 320 && 
b[321] == 321 && 
b[322] == 322 && 
b[323] == 323 && 
b[324] == 324 && 
b[325] == 325 && 
b[326] == 326 && 
b[327] == 327 && 
b[328] == 328 && 
b[329] == 329 && 
b[330] == 330 && 
b[331] == 331 && 
b[332] == 332 && 
b[333] == 333 && 
b[334] == 334 && 
b[335] == 335 && 
b[336] == 336 && 
b[337] == 337 && 
b[338] == 338 && 
b[339] == 339 && 
b[340] == 340 && 
b[341] == 341 && 
b[342] == 342 && 
b[343] == 343 && 
b[344] == 344 && 
b[345] == 345 && 
b[346] == 346 && 
b[347] == 347 && 
b[348] == 348 && 
b[349] == 349 && 
b[350] == 350 && 
b[351] == 351 && 
b[352] == 352 && 
b[353] == 353 && 
b[354] == 354 && 
b[355] == 355 && 
b[356] == 356 && 
b[357] == 357 && 
b[358] == 358 && 
b[359] == 359 && 
b[360] == 360 && 
b[361] == 361 && 
b[362] == 362 && 
b[363] == 363 && 
b[364] == 364 && 
b[365] == 365 && 
b[366] == 366 && 
b[367] == 367 && 
b[368] == 368 && 
b[369] == 369 && 
b[370] == 370 && 
b[371] == 371 && 
b[372] == 372 && 
b[373] == 373 && 
b[374] == 374 && 
b[375] == 375 && 
b[376] == 376 && 
b[377] == 377 && 
b[378] == 378 && 
b[379] == 379 && 
b[380] == 380 && 
b[381] == 381 && 
b[382] == 382 && 
b[383] == 383 && 
b[384] == 384 && 
b[385] == 385 && 
b[386] == 386 && 
b[387] == 387 && 
b[388] == 388 && 
b[389] == 389 && 
b[390] == 390 && 
b[391] == 391 && 
b[392] == 392 && 
b[393] == 393 && 
b[394] == 394 && 
b[395] == 395 && 
b[396] == 396 && 
b[397] == 397 && 
b[398] == 398 && 
b[399] == 399 && 
b[400] == 400 && 
b[401] == 401 && 
b[402] == 402 && 
b[403] == 403 && 
b[404] == 404 && 
b[405] == 405 && 
b[406] == 406 && 
b[407] == 407 && 
b[408] == 408 && 
b[409] == 409 && 
b[410] == 410 && 
b[411] == 411 && 
b[412] == 412 && 
b[413] == 413 && 
b[414] == 414 && 
b[415] == 415 && 
b[416] == 416 && 
b[417] == 417 && 
b[418] == 418 && 
b[419] == 419 && 
b[420] == 420 && 
b[421] == 421 && 
b[422] == 422 && 
b[423] == 423 && 
b[424] == 424 && 
b[425] == 425 && 
b[426] == 426 && 
b[427] == 427 && 
b[428] == 428 && 
b[429] == 429 && 
b[430] == 430 && 
b[431] == 431 && 
b[432] == 432 && 
b[433] == 433 && 
b[434] == 434 && 
b[435] == 435 && 
b[436] == 436 && 
b[437] == 437 && 
b[438] == 438 && 
b[439] == 439 && 
b[440] == 440 && 
b[441] == 441 && 
b[442] == 442 && 
b[443] == 443 && 
b[444] == 444 && 
b[445] == 445 && 
b[446] == 446 && 
b[447] == 447 && 
b[448] == 448 && 
b[449] == 449 && 
b[450] == 450 && 
b[451] == 451 && 
b[452] == 452 && 
b[453] == 453 && 
b[454] == 454 && 
b[455] == 455 && 
b[456] == 456 && 
b[457] == 457 && 
b[458] == 458 && 
b[459] == 459 && 
b[460] == 460 && 
b[461] == 461 && 
b[462] == 462 && 
b[463] == 463 && 
b[464] == 464 && 
b[465] == 465 && 
b[466] == 466 && 
b[467] == 467 && 
b[468] == 468 && 
b[469] == 469 && 
b[470] == 470 && 
b[471] == 471 && 
b[472] == 472 && 
b[473] == 473 && 
b[474] == 474 && 
b[475] == 475 && 
b[476] == 476 && 
b[477] == 477 && 
b[478] == 478 && 
b[479] == 479 && 
b[480] == 480 && 
b[481] == 481 && 
b[482] == 482 && 
b[483] == 483 && 
b[484] == 484 && 
b[485] == 485 && 
b[486] == 486 && 
b[487] == 487 && 
b[488] == 488 && 
b[489] == 489 && 
b[490] == 490 && 
b[491] == 491 && 
b[492] == 492 && 
b[493] == 493 && 
b[494] == 494 && 
b[495] == 495 && 
b[496] == 496 && 
b[497] == 497 && 
b[498] == 498 && 
b[499] == 499 && 
b[500] == 500 && 
b[501] == 501 && 
b[502] == 502 && 
b[503] == 503 && 
b[504] == 504 && 
b[505] == 505 && 
b[506] == 506 && 
b[507] == 507 && 
b[508] == 508 && 
b[509] == 509 && 
b[510] == 510 && 
b[511] == 511 && 
b[512] == 512 && 
b[513] == 513 && 
b[514] == 514 && 
b[515] == 515 && 
b[516] == 516 && 
b[517] == 517 && 
b[518] == 518 && 
b[519] == 519 && 
b[520] == 520 && 
b[521] == 521 && 
b[522] == 522 && 
b[523] == 523 && 
b[524] == 524 && 
b[525] == 525 && 
b[526] == 526 && 
b[527] == 527 && 
b[528] == 528 && 
b[529] == 529 && 
b[530] == 530 && 
b[531] == 531 && 
b[532] == 532 && 
b[533] == 533 && 
b[534] == 534 && 
b[535] == 535 && 
b[536] == 536 && 
b[537] == 537 && 
b[538] == 538 && 
b[539] == 539 && 
b[540] == 540 && 
b[541] == 541 && 
b[542] == 542 && 
b[543] == 543 && 
b[544] == 544 && 
b[545] == 545 && 
b[546] == 546 && 
b[547] == 547 && 
b[548] == 548 && 
b[549] == 549 && 
b[550] == 550 && 
b[551] == 551 && 
b[552] == 552 && 
b[553] == 553 && 
b[554] == 554 && 
b[555] == 555 && 
b[556] == 556 && 
b[557] == 557 && 
b[558] == 558 && 
b[559] == 559 && 
b[560] == 560 && 
b[561] == 561 && 
b[562] == 562 && 
b[563] == 563 && 
b[564] == 564 && 
b[565] == 565 && 
b[566] == 566 && 
b[567] == 567 && 
b[568] == 568 && 
b[569] == 569 && 
b[570] == 570 && 
b[571] == 571 && 
b[572] == 572 && 
b[573] == 573 && 
b[574] == 574 && 
b[575] == 575 && 
b[576] == 576 && 
b[577] == 577 && 
b[578] == 578 && 
b[579] == 579 && 
b[580] == 580 && 
b[581] == 581 && 
b[582] == 582 && 
b[583] == 583 && 
b[584] == 584 && 
b[585] == 585 && 
b[586] == 586 && 
b[587] == 587 && 
b[588] == 588 && 
b[589] == 589 && 
b[590] == 590 && 
b[591] == 591 && 
b[592] == 592 && 
b[593] == 593 && 
b[594] == 594 && 
b[595] == 595 && 
b[596] == 596 && 
b[597] == 597 && 
b[598] == 598 && 
b[599] == 599 && 
b[600] == 600 && 
b[601] == 601 && 
b[602] == 602 && 
b[603] == 603 && 
b[604] == 604 && 
b[605] == 605 && 
b[606] == 606 && 
b[607] == 607 && 
b[608] == 608 && 
b[609] == 609 && 
b[610] == 610 && 
b[611] == 611 && 
b[612] == 612 && 
b[613] == 613 && 
b[614] == 614 && 
b[615] == 615 && 
b[616] == 616 && 
b[617] == 617 && 
b[618] == 618 && 
b[619] == 619 && 
b[620] == 620 && 
b[621] == 621 && 
b[622] == 622 && 
b[623] == 623 && 
b[624] == 624 && 
b[625] == 625 && 
b[626] == 626 && 
b[627] == 627 && 
b[628] == 628 && 
b[629] == 629 && 
b[630] == 630 && 
b[631] == 631 && 
b[632] == 632 && 
b[633] == 633 && 
b[634] == 634 && 
b[635] == 635 && 
b[636] == 636 && 
b[637] == 637 && 
b[638] == 638 && 
b[639] == 639 && 
b[640] == 640 && 
b[641] == 641 && 
b[642] == 642 && 
b[643] == 643 && 
b[644] == 644 && 
b[645] == 645 && 
b[646] == 646 && 
b[647] == 647 && 
b[648] == 648 && 
b[649] == 649 && 
b[650] == 650 && 
b[651] == 651 && 
b[652] == 652 && 
b[653] == 653 && 
b[654] == 654 && 
b[655] == 655 && 
b[656] == 656 && 
b[657] == 657 && 
b[658] == 658 && 
b[659] == 659 && 
b[660] == 660 && 
b[661] == 661 && 
b[662] == 662 && 
b[663] == 663 && 
b[664] == 664 && 
b[665] == 665 && 
b[666] == 666 && 
b[667] == 667 && 
b[668] == 668 && 
b[669] == 669 && 
b[670] == 670 && 
b[671] == 671 && 
b[672] == 672 && 
b[673] == 673 && 
b[674] == 674 && 
b[675] == 675 && 
b[676] == 676 && 
b[677] == 677 && 
b[678] == 678 && 
b[679] == 679 && 
b[680] == 680 && 
b[681] == 681 && 
b[682] == 682 && 
b[683] == 683 && 
b[684] == 684 && 
b[685] == 685 && 
b[686] == 686 && 
b[687] == 687 && 
b[688] == 688 && 
b[689] == 689 && 
b[690] == 690 && 
b[691] == 691 && 
b[692] == 692 && 
b[693] == 693 && 
b[694] == 694 && 
b[695] == 695 && 
b[696] == 696 && 
b[697] == 697 && 
b[698] == 698 && 
b[699] == 699 && 
b[700] == 700 && 
b[701] == 701 && 
b[702] == 702 && 
b[703] == 703 && 
b[704] == 704 && 
b[705] == 705 && 
b[706] == 706 && 
b[707] == 707 && 
b[708] == 708 && 
b[709] == 709 && 
b[710] == 710 && 
b[711] == 711 && 
b[712] == 712 && 
b[713] == 713 && 
b[714] == 714 && 
b[715] == 715 && 
b[716] == 716 && 
b[717] == 717 && 
b[718] == 718 && 
b[719] == 719 && 
b[720] == 720 && 
b[721] == 721 && 
b[722] == 722 && 
b[723] == 723 && 
b[724] == 724 && 
b[725] == 725 && 
b[726] == 726 && 
b[727] == 727 && 
b[728] == 728 && 
b[729] == 729 && 
b[730] == 730 && 
b[731] == 731 && 
b[732] == 732 && 
b[733] == 733 && 
b[734] == 734 && 
b[735] == 735 && 
b[736] == 736 && 
b[737] == 737 && 
b[738] == 738 && 
b[739] == 739 && 
b[740] == 740 && 
b[741] == 741 && 
b[742] == 742 && 
b[743] == 743 && 
b[744] == 744 && 
b[745] == 745 && 
b[746] == 746 && 
b[747] == 747 && 
b[748] == 748 && 
b[749] == 749 && 
b[750] == 750 && 
b[751] == 751 && 
b[752] == 752 && 
b[753] == 753 && 
b[754] == 754 && 
b[755] == 755 && 
b[756] == 756 && 
b[757] == 757 && 
b[758] == 758 && 
b[759] == 759 && 
b[760] == 760 && 
b[761] == 761 && 
b[762] == 762 && 
b[763] == 763 && 
b[764] == 764 && 
b[765] == 765 && 
b[766] == 766 && 
b[767] == 767 && 
b[768] == 768 && 
b[769] == 769 && 
b[770] == 770 && 
b[771] == 771 && 
b[772] == 772 && 
b[773] == 773 && 
b[774] == 774 && 
b[775] == 775 && 
b[776] == 776 && 
b[777] == 777 && 
b[778] == 778 && 
b[779] == 779 && 
b[780] == 780 && 
b[781] == 781 && 
b[782] == 782 && 
b[783] == 783 && 
b[784] == 784 && 
b[785] == 785 && 
b[786] == 786 && 
b[787] == 787 && 
b[788] == 788 && 
b[789] == 789 && 
b[790] == 790 && 
b[791] == 791 && 
b[792] == 792 && 
b[793] == 793 && 
b[794] == 794 && 
b[795] == 795 && 
b[796] == 796 && 
b[797] == 797 && 
b[798] == 798 && 
b[799] == 799 && 
b[800] == 800 && 
b[801] == 801 && 
b[802] == 802 && 
b[803] == 803 && 
b[804] == 804 && 
b[805] == 805 && 
b[806] == 806 && 
b[807] == 807 && 
b[808] == 808 && 
b[809] == 809 && 
b[810] == 810 && 
b[811] == 811 && 
b[812] == 812 && 
b[813] == 813 && 
b[814] == 814 && 
b[815] == 815 && 
b[816] == 816 && 
b[817] == 817 && 
b[818] == 818 && 
b[819] == 819 && 
b[820] == 820 && 
b[821] == 821 && 
b[822] == 822 && 
b[823] == 823 && 
b[824] == 824 && 
b[825] == 825 && 
b[826] == 826 && 
b[827] == 827 && 
b[828] == 828 && 
b[829] == 829 && 
b[830] == 830 && 
b[831] == 831 && 
b[832] == 832 && 
b[833] == 833 && 
b[834] == 834 && 
b[835] == 835 && 
b[836] == 836 && 
b[837] == 837 && 
b[838] == 838 && 
b[839] == 839 && 
b[840] == 840 && 
b[841] == 841 && 
b[842] == 842 && 
b[843] == 843 && 
b[844] == 844 && 
b[845] == 845 && 
b[846] == 846 && 
b[847] == 847 && 
b[848] == 848 && 
b[849] == 849 && 
b[850] == 850 && 
b[851] == 851 && 
b[852] == 852 && 
b[853] == 853 && 
b[854] == 854 && 
b[855] == 855 && 
b[856] == 856 && 
b[857] == 857 && 
b[858] == 858 && 
b[859] == 859 && 
b[860] == 860 && 
b[861] == 861 && 
b[862] == 862 && 
b[863] == 863 && 
b[864] == 864 && 
b[865] == 865 && 
b[866] == 866 && 
b[867] == 867 && 
b[868] == 868 && 
b[869] == 869 && 
b[870] == 870 && 
b[871] == 871 && 
b[872] == 872 && 
b[873] == 873 && 
b[874] == 874 && 
b[875] == 875 && 
b[876] == 876 && 
b[877] == 877 && 
b[878] == 878 && 
b[879] == 879 && 
b[880] == 880 && 
b[881] == 881 && 
b[882] == 882 && 
b[883] == 883 && 
b[884] == 884 && 
b[885] == 885 && 
b[886] == 886 && 
b[887] == 887 && 
b[888] == 888 && 
b[889] == 889 && 
b[890] == 890 && 
b[891] == 891 && 
b[892] == 892 && 
b[893] == 893 && 
b[894] == 894 && 
b[895] == 895 && 
b[896] == 896 && 
b[897] == 897 && 
b[898] == 898 && 
b[899] == 899 && 
b[900] == 900 && 
b[901] == 901 && 
b[902] == 902 && 
b[903] == 903 && 
b[904] == 904 && 
b[905] == 905 && 
b[906] == 906 && 
b[907] == 907 && 
b[908] == 908 && 
b[909] == 909 && 
b[910] == 910 && 
b[911] == 911 && 
b[912] == 912 && 
b[913] == 913 && 
b[914] == 914 && 
b[915] == 915 && 
b[916] == 916 && 
b[917] == 917 && 
b[918] == 918 && 
b[919] == 919 && 
b[920] == 920 && 
b[921] == 921 && 
b[922] == 922 && 
b[923] == 923 && 
b[924] == 924 && 
b[925] == 925 && 
b[926] == 926 && 
b[927] == 927 && 
b[928] == 928 && 
b[929] == 929 && 
b[930] == 930 && 
b[931] == 931 && 
b[932] == 932 && 
b[933] == 933 && 
b[934] == 934 && 
b[935] == 935 && 
b[936] == 936 && 
b[937] == 937 && 
b[938] == 938 && 
b[939] == 939 && 
b[940] == 940 && 
b[941] == 941 && 
b[942] == 942 && 
b[943] == 943 && 
b[944] == 944 && 
b[945] == 945 && 
b[946] == 946 && 
b[947] == 947 && 
b[948] == 948 && 
b[949] == 949 && 
b[950] == 950 && 
b[951] == 951 && 
b[952] == 952 && 
b[953] == 953 && 
b[954] == 954 && 
b[955] == 955 && 
b[956] == 956 && 
b[957] == 957 && 
b[958] == 958 && 
b[959] == 959 && 
b[960] == 960 && 
b[961] == 961 && 
b[962] == 962 && 
b[963] == 963 && 
b[964] == 964 && 
b[965] == 965 && 
b[966] == 966 && 
b[967] == 967 && 
b[968] == 968 && 
b[969] == 969 && 
b[970] == 970 && 
b[971] == 971 && 
b[972] == 972 && 
b[973] == 973 && 
b[974] == 974 && 
b[975] == 975 && 
b[976] == 976 && 
b[977] == 977 && 
b[978] == 978 && 
b[979] == 979 && 
b[980] == 980 && 
b[981] == 981 && 
b[982] == 982 && 
b[983] == 983 && 
b[984] == 984 && 
b[985] == 985 && 
b[986] == 986 && 
b[987] == 987 && 
b[988] == 988 && 
b[989] == 989 && 
b[990] == 990 && 
b[991] == 991 && 
b[992] == 992 && 
b[993] == 993 && 
b[994] == 994 && 
b[995] == 995 && 
b[996] == 996 && 
b[997] == 997 && 
b[998] == 998 && 
b[999] == 999 && 
b[1000] == 1000 && 
b[1001] == 1001 && 
b[1002] == 1002 && 
b[1003] == 1003 && 
b[1004] == 1004 && 
b[1005] == 1005 && 
b[1006] == 1006 && 
b[1007] == 1007 && 
b[1008] == 1008 && 
b[1009] == 1009 && 
b[1010] == 1010 && 
b[1011] == 1011 && 
b[1012] == 1012 && 
b[1013] == 1013 && 
b[1014] == 1014 && 
b[1015] == 1015 && 
b[1016] == 1016 && 
b[1017] == 1017 && 
b[1018] == 1018 && 
b[1019] == 1019 && 
b[1020] == 1020 && 
b[1021] == 1021 && 
b[1022] == 1022 && 
b[1023] == 1023 && 
b[1024] == 1024 && 
b[1025] == 1025 && 
b[1026] == 1026 && 
b[1027] == 1027 && 
b[1028] == 1028 && 
b[1029] == 1029 && 
b[1030] == 1030 && 
b[1031] == 1031 && 
b[1032] == 1032 && 
b[1033] == 1033 && 
b[1034] == 1034 && 
b[1035] == 1035 && 
b[1036] == 1036 && 
b[1037] == 1037 && 
b[1038] == 1038 && 
b[1039] == 1039 && 
b[1040] == 1040 && 
b[1041] == 1041 && 
b[1042] == 1042 && 
b[1043] == 1043 && 
b[1044] == 1044 && 
b[1045] == 1045 && 
b[1046] == 1046 && 
b[1047] == 1047 && 
b[1048] == 1048 && 
b[1049] == 1049 && 
b[1050] == 1050 && 
b[1051] == 1051 && 
b[1052] == 1052 && 
b[1053] == 1053 && 
b[1054] == 1054 && 
b[1055] == 1055 && 
b[1056] == 1056 && 
b[1057] == 1057 && 
b[1058] == 1058 && 
b[1059] == 1059 && 
b[1060] == 1060 && 
b[1061] == 1061 && 
b[1062] == 1062 && 
b[1063] == 1063 && 
b[1064] == 1064 && 
b[1065] == 1065 && 
b[1066] == 1066 && 
b[1067] == 1067 && 
b[1068] == 1068 && 
b[1069] == 1069 && 
b[1070] == 1070 && 
b[1071] == 1071 && 
b[1072] == 1072 && 
b[1073] == 1073 && 
b[1074] == 1074 && 
b[1075] == 1075 && 
b[1076] == 1076 && 
b[1077] == 1077 && 
b[1078] == 1078 && 
b[1079] == 1079 && 
b[1080] == 1080 && 
b[1081] == 1081 && 
b[1082] == 1082 && 
b[1083] == 1083 && 
b[1084] == 1084 && 
b[1085] == 1085 && 
b[1086] == 1086 && 
b[1087] == 1087 && 
b[1088] == 1088 && 
b[1089] == 1089 && 
b[1090] == 1090 && 
b[1091] == 1091 && 
b[1092] == 1092 && 
b[1093] == 1093 && 
b[1094] == 1094 && 
b[1095] == 1095 && 
b[1096] == 1096 && 
b[1097] == 1097 && 
b[1098] == 1098 && 
b[1099] == 1099 && 
b[1100] == 1100 && 
b[1101] == 1101 && 
b[1102] == 1102 && 
b[1103] == 1103 && 
b[1104] == 1104 && 
b[1105] == 1105 && 
b[1106] == 1106 && 
b[1107] == 1107 && 
b[1108] == 1108 && 
b[1109] == 1109 && 
b[1110] == 1110 && 
b[1111] == 1111 && 
b[1112] == 1112 && 
b[1113] == 1113 && 
b[1114] == 1114 && 
b[1115] == 1115 && 
b[1116] == 1116 && 
b[1117] == 1117 && 
b[1118] == 1118 && 
b[1119] == 1119 && 
b[1120] == 1120 && 
b[1121] == 1121 && 
b[1122] == 1122 && 
b[1123] == 1123 && 
b[1124] == 1124 && 
b[1125] == 1125 && 
b[1126] == 1126 && 
b[1127] == 1127 && 
b[1128] == 1128 && 
b[1129] == 1129 && 
b[1130] == 1130 && 
b[1131] == 1131 && 
b[1132] == 1132 && 
b[1133] == 1133 && 
b[1134] == 1134 && 
b[1135] == 1135 && 
b[1136] == 1136 && 
b[1137] == 1137 && 
b[1138] == 1138 && 
b[1139] == 1139 && 
b[1140] == 1140 && 
b[1141] == 1141 && 
b[1142] == 1142 && 
b[1143] == 1143 && 
b[1144] == 1144 && 
b[1145] == 1145 && 
b[1146] == 1146 && 
b[1147] == 1147 && 
b[1148] == 1148 && 
b[1149] == 1149 && 
b[1150] == 1150 && 
b[1151] == 1151 && 
b[1152] == 1152 && 
b[1153] == 1153 && 
b[1154] == 1154 && 
b[1155] == 1155 && 
b[1156] == 1156 && 
b[1157] == 1157 && 
b[1158] == 1158 && 
b[1159] == 1159 && 
b[1160] == 1160 && 
b[1161] == 1161 && 
b[1162] == 1162 && 
b[1163] == 1163 && 
b[1164] == 1164 && 
b[1165] == 1165 && 
b[1166] == 1166 && 
b[1167] == 1167 && 
b[1168] == 1168 && 
b[1169] == 1169 && 
b[1170] == 1170 && 
b[1171] == 1171 && 
b[1172] == 1172 && 
b[1173] == 1173 && 
b[1174] == 1174 && 
b[1175] == 1175 && 
b[1176] == 1176 && 
b[1177] == 1177 && 
b[1178] == 1178 && 
b[1179] == 1179 && 
b[1180] == 1180 && 
b[1181] == 1181 && 
b[1182] == 1182 && 
b[1183] == 1183 && 
b[1184] == 1184 && 
b[1185] == 1185 && 
b[1186] == 1186 && 
b[1187] == 1187 && 
b[1188] == 1188 && 
b[1189] == 1189 && 
b[1190] == 1190 && 
b[1191] == 1191 && 
b[1192] == 1192 && 
b[1193] == 1193 && 
b[1194] == 1194 && 
b[1195] == 1195 && 
b[1196] == 1196 && 
b[1197] == 1197 && 
b[1198] == 1198 && 
b[1199] == 1199 && 
b[1200] == 1200 && 
b[1201] == 1201 && 
b[1202] == 1202 && 
b[1203] == 1203 && 
b[1204] == 1204 && 
b[1205] == 1205 && 
b[1206] == 1206 && 
b[1207] == 1207 && 
b[1208] == 1208 && 
b[1209] == 1209 && 
b[1210] == 1210 && 
b[1211] == 1211 && 
b[1212] == 1212 && 
b[1213] == 1213 && 
b[1214] == 1214 && 
b[1215] == 1215 && 
b[1216] == 1216 && 
b[1217] == 1217 && 
b[1218] == 1218 && 
b[1219] == 1219 && 
b[1220] == 1220 && 
b[1221] == 1221 && 
b[1222] == 1222 && 
b[1223] == 1223 && 
b[1224] == 1224 && 
b[1225] == 1225 && 
b[1226] == 1226 && 
b[1227] == 1227 && 
b[1228] == 1228 && 
b[1229] == 1229 && 
b[1230] == 1230 && 
b[1231] == 1231 && 
b[1232] == 1232 && 
b[1233] == 1233 && 
b[1234] == 1234 && 
b[1235] == 1235 && 
b[1236] == 1236 && 
b[1237] == 1237 && 
b[1238] == 1238 && 
b[1239] == 1239 && 
b[1240] == 1240 && 
b[1241] == 1241 && 
b[1242] == 1242 && 
b[1243] == 1243 && 
b[1244] == 1244 && 
b[1245] == 1245 && 
b[1246] == 1246 && 
b[1247] == 1247 && 
b[1248] == 1248 && 
b[1249] == 1249 && 
b[1250] == 1250 && 
b[1251] == 1251 && 
b[1252] == 1252 && 
b[1253] == 1253 && 
b[1254] == 1254 && 
b[1255] == 1255 && 
b[1256] == 1256 && 
b[1257] == 1257 && 
b[1258] == 1258 && 
b[1259] == 1259 && 
b[1260] == 1260 && 
b[1261] == 1261 && 
b[1262] == 1262 && 
b[1263] == 1263 && 
b[1264] == 1264 && 
b[1265] == 1265 && 
b[1266] == 1266 && 
b[1267] == 1267 && 
b[1268] == 1268 && 
b[1269] == 1269 && 
b[1270] == 1270 && 
b[1271] == 1271 && 
b[1272] == 1272 && 
b[1273] == 1273 && 
b[1274] == 1274 && 
b[1275] == 1275 && 
b[1276] == 1276 && 
b[1277] == 1277 && 
b[1278] == 1278 && 
b[1279] == 1279 && 
b[1280] == 1280 && 
b[1281] == 1281 && 
b[1282] == 1282 && 
b[1283] == 1283 && 
b[1284] == 1284 && 
b[1285] == 1285 && 
b[1286] == 1286 && 
b[1287] == 1287 && 
b[1288] == 1288 && 
b[1289] == 1289 && 
b[1290] == 1290 && 
b[1291] == 1291 && 
b[1292] == 1292 && 
b[1293] == 1293 && 
b[1294] == 1294 && 
b[1295] == 1295 && 
b[1296] == 1296 && 
b[1297] == 1297 && 
b[1298] == 1298 && 
b[1299] == 1299 && 
b[1300] == 1300 && 
b[1301] == 1301 && 
b[1302] == 1302 && 
b[1303] == 1303 && 
b[1304] == 1304 && 
b[1305] == 1305 && 
b[1306] == 1306 && 
b[1307] == 1307 && 
b[1308] == 1308 && 
b[1309] == 1309 && 
b[1310] == 1310 && 
b[1311] == 1311 && 
b[1312] == 1312 && 
b[1313] == 1313 && 
b[1314] == 1314 && 
b[1315] == 1315 && 
b[1316] == 1316 && 
b[1317] == 1317 && 
b[1318] == 1318 && 
b[1319] == 1319 && 
b[1320] == 1320 && 
b[1321] == 1321 && 
b[1322] == 1322 && 
b[1323] == 1323 && 
b[1324] == 1324 && 
b[1325] == 1325 && 
b[1326] == 1326 && 
b[1327] == 1327 && 
b[1328] == 1328 && 
b[1329] == 1329 && 
b[1330] == 1330 && 
b[1331] == 1331 && 
b[1332] == 1332 && 
b[1333] == 1333 && 
b[1334] == 1334 && 
b[1335] == 1335 && 
b[1336] == 1336 && 
b[1337] == 1337 && 
b[1338] == 1338 && 
b[1339] == 1339 && 
b[1340] == 1340 && 
b[1341] == 1341 && 
b[1342] == 1342 && 
b[1343] == 1343 && 
b[1344] == 1344 && 
b[1345] == 1345 && 
b[1346] == 1346 && 
b[1347] == 1347 && 
b[1348] == 1348 && 
b[1349] == 1349 && 
b[1350] == 1350 && 
b[1351] == 1351 && 
b[1352] == 1352 && 
b[1353] == 1353 && 
b[1354] == 1354 && 
b[1355] == 1355 && 
b[1356] == 1356 && 
b[1357] == 1357 && 
b[1358] == 1358 && 
b[1359] == 1359 && 
b[1360] == 1360 && 
b[1361] == 1361 && 
b[1362] == 1362 && 
b[1363] == 1363 && 
b[1364] == 1364 && 
b[1365] == 1365 && 
b[1366] == 1366 && 
b[1367] == 1367 && 
b[1368] == 1368 && 
b[1369] == 1369 && 
b[1370] == 1370 && 
b[1371] == 1371 && 
b[1372] == 1372 && 
b[1373] == 1373 && 
b[1374] == 1374 && 
b[1375] == 1375 && 
b[1376] == 1376 && 
b[1377] == 1377 && 
b[1378] == 1378 && 
b[1379] == 1379 && 
b[1380] == 1380 && 
b[1381] == 1381 && 
b[1382] == 1382 && 
b[1383] == 1383 && 
b[1384] == 1384 && 
b[1385] == 1385 && 
b[1386] == 1386 && 
b[1387] == 1387 && 
b[1388] == 1388 && 
b[1389] == 1389 && 
b[1390] == 1390 && 
b[1391] == 1391 && 
b[1392] == 1392 && 
b[1393] == 1393 && 
b[1394] == 1394 && 
b[1395] == 1395 && 
b[1396] == 1396 && 
b[1397] == 1397 && 
b[1398] == 1398 && 
b[1399] == 1399 && 
b[1400] == 1400 && 
b[1401] == 1401 && 
b[1402] == 1402 && 
b[1403] == 1403 && 
b[1404] == 1404 && 
b[1405] == 1405 && 
b[1406] == 1406 && 
b[1407] == 1407 && 
b[1408] == 1408 && 
b[1409] == 1409 && 
b[1410] == 1410 && 
b[1411] == 1411 && 
b[1412] == 1412 && 
b[1413] == 1413 && 
b[1414] == 1414 && 
b[1415] == 1415 && 
b[1416] == 1416 && 
b[1417] == 1417 && 
b[1418] == 1418 && 
b[1419] == 1419 && 
b[1420] == 1420 && 
b[1421] == 1421 && 
b[1422] == 1422 && 
b[1423] == 1423 && 
b[1424] == 1424 && 
b[1425] == 1425 && 
b[1426] == 1426 && 
b[1427] == 1427 && 
b[1428] == 1428 && 
b[1429] == 1429 && 
b[1430] == 1430 && 
b[1431] == 1431 && 
b[1432] == 1432 && 
b[1433] == 1433 && 
b[1434] == 1434 && 
b[1435] == 1435 && 
b[1436] == 1436 && 
b[1437] == 1437 && 
b[1438] == 1438 && 
b[1439] == 1439 && 
b[1440] == 1440 && 
b[1441] == 1441 && 
b[1442] == 1442 && 
b[1443] == 1443 && 
b[1444] == 1444 && 
b[1445] == 1445 && 
b[1446] == 1446 && 
b[1447] == 1447 && 
b[1448] == 1448 && 
b[1449] == 1449 && 
b[1450] == 1450 && 
b[1451] == 1451 && 
b[1452] == 1452 && 
b[1453] == 1453 && 
b[1454] == 1454 && 
b[1455] == 1455 && 
b[1456] == 1456 && 
b[1457] == 1457 && 
b[1458] == 1458 && 
b[1459] == 1459 && 
b[1460] == 1460 && 
b[1461] == 1461 && 
b[1462] == 1462 && 
b[1463] == 1463 && 
b[1464] == 1464 && 
b[1465] == 1465 && 
b[1466] == 1466 && 
b[1467] == 1467 && 
b[1468] == 1468 && 
b[1469] == 1469 && 
b[1470] == 1470 && 
b[1471] == 1471 && 
b[1472] == 1472 && 
b[1473] == 1473 && 
b[1474] == 1474 && 
b[1475] == 1475 && 
b[1476] == 1476 && 
b[1477] == 1477 && 
b[1478] == 1478 && 
b[1479] == 1479 && 
b[1480] == 1480 && 
b[1481] == 1481 && 
b[1482] == 1482 && 
b[1483] == 1483 && 
b[1484] == 1484 && 
b[1485] == 1485 && 
b[1486] == 1486 && 
b[1487] == 1487 && 
b[1488] == 1488 && 
b[1489] == 1489 && 
b[1490] == 1490 && 
b[1491] == 1491 && 
b[1492] == 1492 && 
b[1493] == 1493 && 
b[1494] == 1494 && 
b[1495] == 1495 && 
b[1496] == 1496 && 
b[1497] == 1497 && 
b[1498] == 1498 && 
b[1499] == 1499 && 
b[1500] == 1500 && 
b[1501] == 1501 && 
b[1502] == 1502 && 
b[1503] == 1503 && 
b[1504] == 1504 && 
b[1505] == 1505 && 
b[1506] == 1506 && 
b[1507] == 1507 && 
b[1508] == 1508 && 
b[1509] == 1509 && 
b[1510] == 1510 && 
b[1511] == 1511 && 
b[1512] == 1512 && 
b[1513] == 1513 && 
b[1514] == 1514 && 
b[1515] == 1515 && 
b[1516] == 1516 && 
b[1517] == 1517 && 
b[1518] == 1518 && 
b[1519] == 1519 && 
b[1520] == 1520 && 
b[1521] == 1521 && 
b[1522] == 1522 && 
b[1523] == 1523 && 
b[1524] == 1524 && 
b[1525] == 1525 && 
b[1526] == 1526 && 
b[1527] == 1527 && 
b[1528] == 1528 && 
b[1529] == 1529 && 
b[1530] == 1530 && 
b[1531] == 1531 && 
b[1532] == 1532 && 
b[1533] == 1533 && 
b[1534] == 1534 && 
b[1535] == 1535 && 
b[1536] == 1536 && 
b[1537] == 1537 && 
b[1538] == 1538 && 
b[1539] == 1539 && 
b[1540] == 1540 && 
b[1541] == 1541 && 
b[1542] == 1542 && 
b[1543] == 1543 && 
b[1544] == 1544 && 
b[1545] == 1545 && 
b[1546] == 1546 && 
b[1547] == 1547 && 
b[1548] == 1548 && 
b[1549] == 1549 && 
b[1550] == 1550 && 
b[1551] == 1551 && 
b[1552] == 1552 && 
b[1553] == 1553 && 
b[1554] == 1554 && 
b[1555] == 1555 && 
b[1556] == 1556 && 
b[1557] == 1557 && 
b[1558] == 1558 && 
b[1559] == 1559 && 
b[1560] == 1560 && 
b[1561] == 1561 && 
b[1562] == 1562 && 
b[1563] == 1563 && 
b[1564] == 1564 && 
b[1565] == 1565 && 
b[1566] == 1566 && 
b[1567] == 1567 && 
b[1568] == 1568 && 
b[1569] == 1569 && 
b[1570] == 1570 && 
b[1571] == 1571 && 
b[1572] == 1572 && 
b[1573] == 1573 && 
b[1574] == 1574 && 
b[1575] == 1575 && 
b[1576] == 1576 && 
b[1577] == 1577 && 
b[1578] == 1578 && 
b[1579] == 1579 && 
b[1580] == 1580 && 
b[1581] == 1581 && 
b[1582] == 1582 && 
b[1583] == 1583 && 
b[1584] == 1584 && 
b[1585] == 1585 && 
b[1586] == 1586 && 
b[1587] == 1587 && 
b[1588] == 1588 && 
b[1589] == 1589 && 
b[1590] == 1590 && 
b[1591] == 1591 && 
b[1592] == 1592 && 
b[1593] == 1593 && 
b[1594] == 1594 && 
b[1595] == 1595 && 
b[1596] == 1596 && 
b[1597] == 1597 && 
b[1598] == 1598 && 
b[1599] == 1599 && 
b[1600] == 1600 && 
b[1601] == 1601 && 
b[1602] == 1602 && 
b[1603] == 1603 && 
b[1604] == 1604 && 
b[1605] == 1605 && 
b[1606] == 1606 && 
b[1607] == 1607 && 
b[1608] == 1608 && 
b[1609] == 1609 && 
b[1610] == 1610 && 
b[1611] == 1611 && 
b[1612] == 1612 && 
b[1613] == 1613 && 
b[1614] == 1614 && 
b[1615] == 1615 && 
b[1616] == 1616 && 
b[1617] == 1617 && 
b[1618] == 1618 && 
b[1619] == 1619 && 
b[1620] == 1620 && 
b[1621] == 1621 && 
b[1622] == 1622 && 
b[1623] == 1623 && 
b[1624] == 1624 && 
b[1625] == 1625 && 
b[1626] == 1626 && 
b[1627] == 1627 && 
b[1628] == 1628 && 
b[1629] == 1629 && 
b[1630] == 1630 && 
b[1631] == 1631 && 
b[1632] == 1632 && 
b[1633] == 1633 && 
b[1634] == 1634 && 
b[1635] == 1635 && 
b[1636] == 1636 && 
b[1637] == 1637 && 
b[1638] == 1638 && 
b[1639] == 1639 && 
b[1640] == 1640 && 
b[1641] == 1641 && 
b[1642] == 1642 && 
b[1643] == 1643 && 
b[1644] == 1644 && 
b[1645] == 1645 && 
b[1646] == 1646 && 
b[1647] == 1647 && 
b[1648] == 1648 && 
b[1649] == 1649 && 
b[1650] == 1650 && 
b[1651] == 1651 && 
b[1652] == 1652 && 
b[1653] == 1653 && 
b[1654] == 1654 && 
b[1655] == 1655 && 
b[1656] == 1656 && 
b[1657] == 1657 && 
b[1658] == 1658 && 
b[1659] == 1659 && 
b[1660] == 1660 && 
b[1661] == 1661 && 
b[1662] == 1662 && 
b[1663] == 1663 && 
b[1664] == 1664 && 
b[1665] == 1665 && 
b[1666] == 1666 && 
b[1667] == 1667 && 
b[1668] == 1668 && 
b[1669] == 1669 && 
b[1670] == 1670 && 
b[1671] == 1671 && 
b[1672] == 1672 && 
b[1673] == 1673 && 
b[1674] == 1674 && 
b[1675] == 1675 && 
b[1676] == 1676 && 
b[1677] == 1677 && 
b[1678] == 1678 && 
b[1679] == 1679 && 
b[1680] == 1680 && 
b[1681] == 1681 && 
b[1682] == 1682 && 
b[1683] == 1683 && 
b[1684] == 1684 && 
b[1685] == 1685 && 
b[1686] == 1686 && 
b[1687] == 1687 && 
b[1688] == 1688 && 
b[1689] == 1689 && 
b[1690] == 1690 && 
b[1691] == 1691 && 
b[1692] == 1692 && 
b[1693] == 1693 && 
b[1694] == 1694 && 
b[1695] == 1695 && 
b[1696] == 1696 && 
b[1697] == 1697 && 
b[1698] == 1698 && 
b[1699] == 1699 && 
b[1700] == 1700 && 
b[1701] == 1701 && 
b[1702] == 1702 && 
b[1703] == 1703 && 
b[1704] == 1704 && 
b[1705] == 1705 && 
b[1706] == 1706 && 
b[1707] == 1707 && 
b[1708] == 1708 && 
b[1709] == 1709 && 
b[1710] == 1710 && 
b[1711] == 1711 && 
b[1712] == 1712 && 
b[1713] == 1713 && 
b[1714] == 1714 && 
b[1715] == 1715 && 
b[1716] == 1716 && 
b[1717] == 1717 && 
b[1718] == 1718 && 
b[1719] == 1719 && 
b[1720] == 1720 && 
b[1721] == 1721 && 
b[1722] == 1722 && 
b[1723] == 1723 && 
b[1724] == 1724 && 
b[1725] == 1725 && 
b[1726] == 1726 && 
b[1727] == 1727 && 
b[1728] == 1728 && 
b[1729] == 1729 && 
b[1730] == 1730 && 
b[1731] == 1731 && 
b[1732] == 1732 && 
b[1733] == 1733 && 
b[1734] == 1734 && 
b[1735] == 1735 && 
b[1736] == 1736 && 
b[1737] == 1737 && 
b[1738] == 1738 && 
b[1739] == 1739 && 
b[1740] == 1740 && 
b[1741] == 1741 && 
b[1742] == 1742 && 
b[1743] == 1743 && 
b[1744] == 1744 && 
b[1745] == 1745 && 
b[1746] == 1746 && 
b[1747] == 1747 && 
b[1748] == 1748 && 
b[1749] == 1749 && 
b[1750] == 1750 && 
b[1751] == 1751 && 
b[1752] == 1752 && 
b[1753] == 1753 && 
b[1754] == 1754 && 
b[1755] == 1755 && 
b[1756] == 1756 && 
b[1757] == 1757 && 
b[1758] == 1758 && 
b[1759] == 1759 && 
b[1760] == 1760 && 
b[1761] == 1761 && 
b[1762] == 1762 && 
b[1763] == 1763 && 
b[1764] == 1764 && 
b[1765] == 1765 && 
b[1766] == 1766 && 
b[1767] == 1767 && 
b[1768] == 1768 && 
b[1769] == 1769 && 
b[1770] == 1770 && 
b[1771] == 1771 && 
b[1772] == 1772 && 
b[1773] == 1773 && 
b[1774] == 1774 && 
b[1775] == 1775 && 
b[1776] == 1776 && 
b[1777] == 1777 && 
b[1778] == 1778 && 
b[1779] == 1779 && 
b[1780] == 1780 && 
b[1781] == 1781 && 
b[1782] == 1782 && 
b[1783] == 1783 && 
b[1784] == 1784 && 
b[1785] == 1785 && 
b[1786] == 1786 && 
b[1787] == 1787 && 
b[1788] == 1788 && 
b[1789] == 1789 && 
b[1790] == 1790 && 
b[1791] == 1791 && 
b[1792] == 1792 && 
b[1793] == 1793 && 
b[1794] == 1794 && 
b[1795] == 1795 && 
b[1796] == 1796 && 
b[1797] == 1797 && 
b[1798] == 1798 && 
b[1799] == 1799 && 
b[1800] == 1800 && 
b[1801] == 1801 && 
b[1802] == 1802 && 
b[1803] == 1803 && 
b[1804] == 1804 && 
b[1805] == 1805 && 
b[1806] == 1806 && 
b[1807] == 1807 && 
b[1808] == 1808 && 
b[1809] == 1809 && 
b[1810] == 1810 && 
b[1811] == 1811 && 
b[1812] == 1812 && 
b[1813] == 1813 && 
b[1814] == 1814 && 
b[1815] == 1815 && 
b[1816] == 1816 && 
b[1817] == 1817 && 
b[1818] == 1818 && 
b[1819] == 1819 && 
b[1820] == 1820 && 
b[1821] == 1821 && 
b[1822] == 1822 && 
b[1823] == 1823 && 
b[1824] == 1824 && 
b[1825] == 1825 && 
b[1826] == 1826 && 
b[1827] == 1827 && 
b[1828] == 1828 && 
b[1829] == 1829 && 
b[1830] == 1830 && 
b[1831] == 1831 && 
b[1832] == 1832 && 
b[1833] == 1833 && 
b[1834] == 1834 && 
b[1835] == 1835 && 
b[1836] == 1836 && 
b[1837] == 1837 && 
b[1838] == 1838 && 
b[1839] == 1839 && 
b[1840] == 1840 && 
b[1841] == 1841 && 
b[1842] == 1842 && 
b[1843] == 1843 && 
b[1844] == 1844 && 
b[1845] == 1845 && 
b[1846] == 1846 && 
b[1847] == 1847 && 
b[1848] == 1848 && 
b[1849] == 1849 && 
b[1850] == 1850 && 
b[1851] == 1851 && 
b[1852] == 1852 && 
b[1853] == 1853 && 
b[1854] == 1854 && 
b[1855] == 1855 && 
b[1856] == 1856 && 
b[1857] == 1857 && 
b[1858] == 1858 && 
b[1859] == 1859 && 
b[1860] == 1860 && 
b[1861] == 1861 && 
b[1862] == 1862 && 
b[1863] == 1863 && 
b[1864] == 1864 && 
b[1865] == 1865 && 
b[1866] == 1866 && 
b[1867] == 1867 && 
b[1868] == 1868 && 
b[1869] == 1869 && 
b[1870] == 1870 && 
b[1871] == 1871 && 
b[1872] == 1872 && 
b[1873] == 1873 && 
b[1874] == 1874 && 
b[1875] == 1875 && 
b[1876] == 1876 && 
b[1877] == 1877 && 
b[1878] == 1878 && 
b[1879] == 1879 && 
b[1880] == 1880 && 
b[1881] == 1881 && 
b[1882] == 1882 && 
b[1883] == 1883 && 
b[1884] == 1884 && 
b[1885] == 1885 && 
b[1886] == 1886 && 
b[1887] == 1887 && 
b[1888] == 1888 && 
b[1889] == 1889 && 
b[1890] == 1890 && 
b[1891] == 1891 && 
b[1892] == 1892 && 
b[1893] == 1893 && 
b[1894] == 1894 && 
b[1895] == 1895 && 
b[1896] == 1896 && 
b[1897] == 1897 && 
b[1898] == 1898 && 
b[1899] == 1899 && 
b[1900] == 1900 && 
b[1901] == 1901 && 
b[1902] == 1902 && 
b[1903] == 1903 && 
b[1904] == 1904 && 
b[1905] == 1905 && 
b[1906] == 1906 && 
b[1907] == 1907 && 
b[1908] == 1908 && 
b[1909] == 1909 && 
b[1910] == 1910 && 
b[1911] == 1911 && 
b[1912] == 1912 && 
b[1913] == 1913 && 
b[1914] == 1914 && 
b[1915] == 1915 && 
b[1916] == 1916 && 
b[1917] == 1917 && 
b[1918] == 1918 && 
b[1919] == 1919 && 
b[1920] == 1920 && 
b[1921] == 1921 && 
b[1922] == 1922 && 
b[1923] == 1923 && 
b[1924] == 1924 && 
b[1925] == 1925 && 
b[1926] == 1926 && 
b[1927] == 1927 && 
b[1928] == 1928 && 
b[1929] == 1929 && 
b[1930] == 1930 && 
b[1931] == 1931 && 
b[1932] == 1932 && 
b[1933] == 1933 && 
b[1934] == 1934 && 
b[1935] == 1935 && 
b[1936] == 1936 && 
b[1937] == 1937 && 
b[1938] == 1938 && 
b[1939] == 1939 && 
b[1940] == 1940 && 
b[1941] == 1941 && 
b[1942] == 1942 && 
b[1943] == 1943 && 
b[1944] == 1944 && 
b[1945] == 1945 && 
b[1946] == 1946 && 
b[1947] == 1947 && 
b[1948] == 1948 && 
b[1949] == 1949 && 
b[1950] == 1950 && 
b[1951] == 1951 && 
b[1952] == 1952 && 
b[1953] == 1953 && 
b[1954] == 1954 && 
b[1955] == 1955 && 
b[1956] == 1956 && 
b[1957] == 1957 && 
b[1958] == 1958 && 
b[1959] == 1959 && 
b[1960] == 1960 && 
b[1961] == 1961 && 
b[1962] == 1962 && 
b[1963] == 1963 && 
b[1964] == 1964 && 
b[1965] == 1965 && 
b[1966] == 1966 && 
b[1967] == 1967 && 
b[1968] == 1968 && 
b[1969] == 1969 && 
b[1970] == 1970 && 
b[1971] == 1971 && 
b[1972] == 1972 && 
b[1973] == 1973 && 
b[1974] == 1974 && 
b[1975] == 1975 && 
b[1976] == 1976 && 
b[1977] == 1977 && 
b[1978] == 1978 && 
b[1979] == 1979 && 
b[1980] == 1980 && 
b[1981] == 1981 && 
b[1982] == 1982 && 
b[1983] == 1983 && 
b[1984] == 1984 && 
b[1985] == 1985 && 
b[1986] == 1986 && 
b[1987] == 1987 && 
b[1988] == 1988 && 
b[1989] == 1989 && 
b[1990] == 1990 && 
b[1991] == 1991 && 
b[1992] == 1992 && 
b[1993] == 1993 && 
b[1994] == 1994 && 
b[1995] == 1995 && 
b[1996] == 1996 && 
b[1997] == 1997 && 
b[1998] == 1998 && 
b[1999] == 1999 && 
b[2000] == 2000 && 
b[2001] == 2001 && 
b[2002] == 2002 && 
b[2003] == 2003 && 
b[2004] == 2004 && 
b[2005] == 2005 && 
b[2006] == 2006 && 
b[2007] == 2007 && 
b[2008] == 2008 && 
b[2009] == 2009 && 
b[2010] == 2010 && 
b[2011] == 2011 && 
b[2012] == 2012 && 
b[2013] == 2013 && 
b[2014] == 2014 && 
b[2015] == 2015 && 
b[2016] == 2016 && 
b[2017] == 2017 && 
b[2018] == 2018 && 
b[2019] == 2019 && 
b[2020] == 2020 && 
b[2021] == 2021 && 
b[2022] == 2022 && 
b[2023] == 2023 && 
b[2024] == 2024 && 
b[2025] == 2025 && 
b[2026] == 2026 && 
b[2027] == 2027 && 
b[2028] == 2028 && 
b[2029] == 2029 && 
b[2030] == 2030 && 
b[2031] == 2031 && 
b[2032] == 2032 && 
b[2033] == 2033 && 
b[2034] == 2034 && 
b[2035] == 2035 && 
b[2036] == 2036 && 
b[2037] == 2037 && 
b[2038] == 2038 && 
b[2039] == 2039 && 
b[2040] == 2040 && 
b[2041] == 2041 && 
b[2042] == 2042 && 
b[2043] == 2043 && 
b[2044] == 2044 && 
b[2045] == 2045 && 
b[2046] == 2046 && 
b[2047] == 2047 && 
b[2048] == 2048 && 
b[2049] == 2049 && 
b[2050] == 2050 && 
b[2051] == 2051 && 
b[2052] == 2052 && 
b[2053] == 2053 && 
b[2054] == 2054 && 
b[2055] == 2055 && 
b[2056] == 2056 && 
b[2057] == 2057 && 
b[2058] == 2058 && 
b[2059] == 2059 && 
b[2060] == 2060 && 
b[2061] == 2061 && 
b[2062] == 2062 && 
b[2063] == 2063 && 
b[2064] == 2064 && 
b[2065] == 2065 && 
b[2066] == 2066 && 
b[2067] == 2067 && 
b[2068] == 2068 && 
b[2069] == 2069 && 
b[2070] == 2070 && 
b[2071] == 2071 && 
b[2072] == 2072 && 
b[2073] == 2073 && 
b[2074] == 2074 && 
b[2075] == 2075 && 
b[2076] == 2076 && 
b[2077] == 2077 && 
b[2078] == 2078 && 
b[2079] == 2079 && 
b[2080] == 2080 && 
b[2081] == 2081 && 
b[2082] == 2082 && 
b[2083] == 2083 && 
b[2084] == 2084 && 
b[2085] == 2085 && 
b[2086] == 2086 && 
b[2087] == 2087 && 
b[2088] == 2088 && 
b[2089] == 2089 && 
b[2090] == 2090 && 
b[2091] == 2091 && 
b[2092] == 2092 && 
b[2093] == 2093 && 
b[2094] == 2094 && 
b[2095] == 2095 && 
b[2096] == 2096 && 
b[2097] == 2097 && 
b[2098] == 2098 && 
b[2099] == 2099 && 
b[2100] == 2100 && 
b[2101] == 2101 && 
b[2102] == 2102 && 
b[2103] == 2103 && 
b[2104] == 2104 && 
b[2105] == 2105 && 
b[2106] == 2106 && 
b[2107] == 2107 && 
b[2108] == 2108 && 
b[2109] == 2109 && 
b[2110] == 2110 && 
b[2111] == 2111 && 
b[2112] == 2112 && 
b[2113] == 2113 && 
b[2114] == 2114 && 
b[2115] == 2115 && 
b[2116] == 2116 && 
b[2117] == 2117 && 
b[2118] == 2118 && 
b[2119] == 2119 && 
b[2120] == 2120 && 
b[2121] == 2121 && 
b[2122] == 2122 && 
b[2123] == 2123 && 
b[2124] == 2124 && 
b[2125] == 2125 && 
b[2126] == 2126 && 
b[2127] == 2127 && 
b[2128] == 2128 && 
b[2129] == 2129 && 
b[2130] == 2130 && 
b[2131] == 2131 && 
b[2132] == 2132 && 
b[2133] == 2133 && 
b[2134] == 2134 && 
b[2135] == 2135 && 
b[2136] == 2136 && 
b[2137] == 2137 && 
b[2138] == 2138 && 
b[2139] == 2139 && 
b[2140] == 2140 && 
b[2141] == 2141 && 
b[2142] == 2142 && 
b[2143] == 2143 && 
b[2144] == 2144 && 
b[2145] == 2145 && 
b[2146] == 2146 && 
b[2147] == 2147 && 
b[2148] == 2148 && 
b[2149] == 2149 && 
b[2150] == 2150 && 
b[2151] == 2151 && 
b[2152] == 2152 && 
b[2153] == 2153 && 
b[2154] == 2154 && 
b[2155] == 2155 && 
b[2156] == 2156 && 
b[2157] == 2157 && 
b[2158] == 2158 && 
b[2159] == 2159 && 
b[2160] == 2160 && 
b[2161] == 2161 && 
b[2162] == 2162 && 
b[2163] == 2163 && 
b[2164] == 2164 && 
b[2165] == 2165 && 
b[2166] == 2166 && 
b[2167] == 2167 && 
b[2168] == 2168 && 
b[2169] == 2169 && 
b[2170] == 2170 && 
b[2171] == 2171 && 
b[2172] == 2172 && 
b[2173] == 2173 && 
b[2174] == 2174 && 
b[2175] == 2175 && 
b[2176] == 2176 && 
b[2177] == 2177 && 
b[2178] == 2178 && 
b[2179] == 2179 && 
b[2180] == 2180 && 
b[2181] == 2181 && 
b[2182] == 2182 && 
b[2183] == 2183 && 
b[2184] == 2184 && 
b[2185] == 2185 && 
b[2186] == 2186 && 
b[2187] == 2187 && 
b[2188] == 2188 && 
b[2189] == 2189 && 
b[2190] == 2190 && 
b[2191] == 2191 && 
b[2192] == 2192 && 
b[2193] == 2193 && 
b[2194] == 2194 && 
b[2195] == 2195 && 
b[2196] == 2196 && 
b[2197] == 2197 && 
b[2198] == 2198 && 
b[2199] == 2199 && 
b[2200] == 2200 && 
b[2201] == 2201 && 
b[2202] == 2202 && 
b[2203] == 2203 && 
b[2204] == 2204 && 
b[2205] == 2205 && 
b[2206] == 2206 && 
b[2207] == 2207 && 
b[2208] == 2208 && 
b[2209] == 2209 && 
b[2210] == 2210 && 
b[2211] == 2211 && 
b[2212] == 2212 && 
b[2213] == 2213 && 
b[2214] == 2214 && 
b[2215] == 2215 && 
b[2216] == 2216 && 
b[2217] == 2217 && 
b[2218] == 2218 && 
b[2219] == 2219 && 
b[2220] == 2220 && 
b[2221] == 2221 && 
b[2222] == 2222 && 
b[2223] == 2223 && 
b[2224] == 2224 && 
b[2225] == 2225 && 
b[2226] == 2226 && 
b[2227] == 2227 && 
b[2228] == 2228 && 
b[2229] == 2229 && 
b[2230] == 2230 && 
b[2231] == 2231 && 
b[2232] == 2232 && 
b[2233] == 2233 && 
b[2234] == 2234 && 
b[2235] == 2235 && 
b[2236] == 2236 && 
b[2237] == 2237 && 
b[2238] == 2238 && 
b[2239] == 2239 && 
b[2240] == 2240 && 
b[2241] == 2241 && 
b[2242] == 2242 && 
b[2243] == 2243 && 
b[2244] == 2244 && 
b[2245] == 2245 && 
b[2246] == 2246 && 
b[2247] == 2247 && 
b[2248] == 2248 && 
b[2249] == 2249 && 
b[2250] == 2250 && 
b[2251] == 2251 && 
b[2252] == 2252 && 
b[2253] == 2253 && 
b[2254] == 2254 && 
b[2255] == 2255 && 
b[2256] == 2256 && 
b[2257] == 2257 && 
b[2258] == 2258 && 
b[2259] == 2259 && 
b[2260] == 2260 && 
b[2261] == 2261 && 
b[2262] == 2262 && 
b[2263] == 2263 && 
b[2264] == 2264 && 
b[2265] == 2265 && 
b[2266] == 2266 && 
b[2267] == 2267 && 
b[2268] == 2268 && 
b[2269] == 2269 && 
b[2270] == 2270 && 
b[2271] == 2271 && 
b[2272] == 2272 && 
b[2273] == 2273 && 
b[2274] == 2274 && 
b[2275] == 2275 && 
b[2276] == 2276 && 
b[2277] == 2277 && 
b[2278] == 2278 && 
b[2279] == 2279 && 
b[2280] == 2280 && 
b[2281] == 2281 && 
b[2282] == 2282 && 
b[2283] == 2283 && 
b[2284] == 2284 && 
b[2285] == 2285 && 
b[2286] == 2286 && 
b[2287] == 2287 && 
b[2288] == 2288 && 
b[2289] == 2289 && 
b[2290] == 2290 && 
b[2291] == 2291 && 
b[2292] == 2292 && 
b[2293] == 2293 && 
b[2294] == 2294 && 
b[2295] == 2295 && 
b[2296] == 2296 && 
b[2297] == 2297 && 
b[2298] == 2298 && 
b[2299] == 2299 && 
b[2300] == 2300 && 
b[2301] == 2301 && 
b[2302] == 2302 && 
b[2303] == 2303 && 
b[2304] == 2304 && 
b[2305] == 2305 && 
b[2306] == 2306 && 
b[2307] == 2307 && 
b[2308] == 2308 && 
b[2309] == 2309 && 
b[2310] == 2310 && 
b[2311] == 2311 && 
b[2312] == 2312 && 
b[2313] == 2313 && 
b[2314] == 2314 && 
b[2315] == 2315 && 
b[2316] == 2316 && 
b[2317] == 2317 && 
b[2318] == 2318 && 
b[2319] == 2319 && 
b[2320] == 2320 && 
b[2321] == 2321 && 
b[2322] == 2322 && 
b[2323] == 2323 && 
b[2324] == 2324 && 
b[2325] == 2325 && 
b[2326] == 2326 && 
b[2327] == 2327 && 
b[2328] == 2328 && 
b[2329] == 2329 && 
b[2330] == 2330 && 
b[2331] == 2331 && 
b[2332] == 2332 && 
b[2333] == 2333 && 
b[2334] == 2334 && 
b[2335] == 2335 && 
b[2336] == 2336 && 
b[2337] == 2337 && 
b[2338] == 2338 && 
b[2339] == 2339 && 
b[2340] == 2340 && 
b[2341] == 2341 && 
b[2342] == 2342 && 
b[2343] == 2343 && 
b[2344] == 2344 && 
b[2345] == 2345 && 
b[2346] == 2346 && 
b[2347] == 2347 && 
b[2348] == 2348 && 
b[2349] == 2349 && 
b[2350] == 2350 && 
b[2351] == 2351 && 
b[2352] == 2352 && 
b[2353] == 2353 && 
b[2354] == 2354 && 
b[2355] == 2355 && 
b[2356] == 2356 && 
b[2357] == 2357 && 
b[2358] == 2358 && 
b[2359] == 2359 && 
b[2360] == 2360 && 
b[2361] == 2361 && 
b[2362] == 2362 && 
b[2363] == 2363 && 
b[2364] == 2364 && 
b[2365] == 2365 && 
b[2366] == 2366 && 
b[2367] == 2367 && 
b[2368] == 2368 && 
b[2369] == 2369 && 
b[2370] == 2370 && 
b[2371] == 2371 && 
b[2372] == 2372 && 
b[2373] == 2373 && 
b[2374] == 2374 && 
b[2375] == 2375 && 
b[2376] == 2376 && 
b[2377] == 2377 && 
b[2378] == 2378 && 
b[2379] == 2379 && 
b[2380] == 2380 && 
b[2381] == 2381 && 
b[2382] == 2382 && 
b[2383] == 2383 && 
b[2384] == 2384 && 
b[2385] == 2385 && 
b[2386] == 2386 && 
b[2387] == 2387 && 
b[2388] == 2388 && 
b[2389] == 2389 && 
b[2390] == 2390 && 
b[2391] == 2391 && 
b[2392] == 2392 && 
b[2393] == 2393 && 
b[2394] == 2394 && 
b[2395] == 2395 && 
b[2396] == 2396 && 
b[2397] == 2397 && 
b[2398] == 2398 && 
b[2399] == 2399 && 
b[2400] == 2400 && 
b[2401] == 2401 && 
b[2402] == 2402 && 
b[2403] == 2403 && 
b[2404] == 2404 && 
b[2405] == 2405 && 
b[2406] == 2406 && 
b[2407] == 2407 && 
b[2408] == 2408 && 
b[2409] == 2409 && 
b[2410] == 2410 && 
b[2411] == 2411 && 
b[2412] == 2412 && 
b[2413] == 2413 && 
b[2414] == 2414 && 
b[2415] == 2415 && 
b[2416] == 2416 && 
b[2417] == 2417 && 
b[2418] == 2418 && 
b[2419] == 2419 && 
b[2420] == 2420 && 
b[2421] == 2421 && 
b[2422] == 2422 && 
b[2423] == 2423 && 
b[2424] == 2424 && 
b[2425] == 2425 && 
b[2426] == 2426 && 
b[2427] == 2427 && 
b[2428] == 2428 && 
b[2429] == 2429 && 
b[2430] == 2430 && 
b[2431] == 2431 && 
b[2432] == 2432 && 
b[2433] == 2433 && 
b[2434] == 2434 && 
b[2435] == 2435 && 
b[2436] == 2436 && 
b[2437] == 2437 && 
b[2438] == 2438 && 
b[2439] == 2439 && 
b[2440] == 2440 && 
b[2441] == 2441 && 
b[2442] == 2442 && 
b[2443] == 2443 && 
b[2444] == 2444 && 
b[2445] == 2445 && 
b[2446] == 2446 && 
b[2447] == 2447 && 
b[2448] == 2448 && 
b[2449] == 2449 && 
b[2450] == 2450 && 
b[2451] == 2451 && 
b[2452] == 2452 && 
b[2453] == 2453 && 
b[2454] == 2454 && 
b[2455] == 2455 && 
b[2456] == 2456 && 
b[2457] == 2457 && 
b[2458] == 2458 && 
b[2459] == 2459 && 
b[2460] == 2460 && 
b[2461] == 2461 && 
b[2462] == 2462 && 
b[2463] == 2463 && 
b[2464] == 2464 && 
b[2465] == 2465 && 
b[2466] == 2466 && 
b[2467] == 2467 && 
b[2468] == 2468 && 
b[2469] == 2469 && 
b[2470] == 2470 && 
b[2471] == 2471 && 
b[2472] == 2472 && 
b[2473] == 2473 && 
b[2474] == 2474 && 
b[2475] == 2475 && 
b[2476] == 2476 && 
b[2477] == 2477 && 
b[2478] == 2478 && 
b[2479] == 2479 && 
b[2480] == 2480 && 
b[2481] == 2481 && 
b[2482] == 2482 && 
b[2483] == 2483 && 
b[2484] == 2484 && 
b[2485] == 2485 && 
b[2486] == 2486 && 
b[2487] == 2487 && 
b[2488] == 2488 && 
b[2489] == 2489 && 
b[2490] == 2490 && 
b[2491] == 2491 && 
b[2492] == 2492 && 
b[2493] == 2493 && 
b[2494] == 2494 && 
b[2495] == 2495 && 
b[2496] == 2496 && 
b[2497] == 2497 && 
b[2498] == 2498 && 
b[2499] == 2499 && 
b[2500] == 2500 && 
b[2501] == 2501 && 
b[2502] == 2502 && 
b[2503] == 2503 && 
b[2504] == 2504 && 
b[2505] == 2505 && 
b[2506] == 2506 && 
b[2507] == 2507 && 
b[2508] == 2508 && 
b[2509] == 2509 && 
b[2510] == 2510 && 
b[2511] == 2511 && 
b[2512] == 2512 && 
b[2513] == 2513 && 
b[2514] == 2514 && 
b[2515] == 2515 && 
b[2516] == 2516 && 
b[2517] == 2517 && 
b[2518] == 2518 && 
b[2519] == 2519 && 
b[2520] == 2520 && 
b[2521] == 2521 && 
b[2522] == 2522 && 
b[2523] == 2523 && 
b[2524] == 2524 && 
b[2525] == 2525 && 
b[2526] == 2526 && 
b[2527] == 2527 && 
b[2528] == 2528 && 
b[2529] == 2529 && 
b[2530] == 2530 && 
b[2531] == 2531 && 
b[2532] == 2532 && 
b[2533] == 2533 && 
b[2534] == 2534 && 
b[2535] == 2535 && 
b[2536] == 2536 && 
b[2537] == 2537 && 
b[2538] == 2538 && 
b[2539] == 2539 && 
b[2540] == 2540 && 
b[2541] == 2541 && 
b[2542] == 2542 && 
b[2543] == 2543 && 
b[2544] == 2544 && 
b[2545] == 2545 && 
b[2546] == 2546 && 
b[2547] == 2547 && 
b[2548] == 2548 && 
b[2549] == 2549 && 
b[2550] == 2550 && 
b[2551] == 2551 && 
b[2552] == 2552 && 
b[2553] == 2553 && 
b[2554] == 2554 && 
b[2555] == 2555 && 
b[2556] == 2556 && 
b[2557] == 2557 && 
b[2558] == 2558 && 
b[2559] == 2559 && 
b[2560] == 2560 && 
b[2561] == 2561 && 
b[2562] == 2562 && 
b[2563] == 2563 && 
b[2564] == 2564 && 
b[2565] == 2565 && 
b[2566] == 2566 && 
b[2567] == 2567 && 
b[2568] == 2568 && 
b[2569] == 2569 && 
b[2570] == 2570 && 
b[2571] == 2571 && 
b[2572] == 2572 && 
b[2573] == 2573 && 
b[2574] == 2574 && 
b[2575] == 2575 && 
b[2576] == 2576 && 
b[2577] == 2577 && 
b[2578] == 2578 && 
b[2579] == 2579 && 
b[2580] == 2580 && 
b[2581] == 2581 && 
b[2582] == 2582 && 
b[2583] == 2583 && 
b[2584] == 2584 && 
b[2585] == 2585 && 
b[2586] == 2586 && 
b[2587] == 2587 && 
b[2588] == 2588 && 
b[2589] == 2589 && 
b[2590] == 2590 && 
b[2591] == 2591 && 
b[2592] == 2592 && 
b[2593] == 2593 && 
b[2594] == 2594 && 
b[2595] == 2595 && 
b[2596] == 2596 && 
b[2597] == 2597 && 
b[2598] == 2598 && 
b[2599] == 2599 && 
b[2600] == 2600 && 
b[2601] == 2601 && 
b[2602] == 2602 && 
b[2603] == 2603 && 
b[2604] == 2604 && 
b[2605] == 2605 && 
b[2606] == 2606 && 
b[2607] == 2607 && 
b[2608] == 2608 && 
b[2609] == 2609 && 
b[2610] == 2610 && 
b[2611] == 2611 && 
b[2612] == 2612 && 
b[2613] == 2613 && 
b[2614] == 2614 && 
b[2615] == 2615 && 
b[2616] == 2616 && 
b[2617] == 2617 && 
b[2618] == 2618 && 
b[2619] == 2619 && 
b[2620] == 2620 && 
b[2621] == 2621 && 
b[2622] == 2622 && 
b[2623] == 2623 && 
b[2624] == 2624 && 
b[2625] == 2625 && 
b[2626] == 2626 && 
b[2627] == 2627 && 
b[2628] == 2628 && 
b[2629] == 2629 && 
b[2630] == 2630 && 
b[2631] == 2631 && 
b[2632] == 2632 && 
b[2633] == 2633 && 
b[2634] == 2634 && 
b[2635] == 2635 && 
b[2636] == 2636 && 
b[2637] == 2637 && 
b[2638] == 2638 && 
b[2639] == 2639 && 
b[2640] == 2640 && 
b[2641] == 2641 && 
b[2642] == 2642 && 
b[2643] == 2643 && 
b[2644] == 2644 && 
b[2645] == 2645 && 
b[2646] == 2646 && 
b[2647] == 2647 && 
b[2648] == 2648 && 
b[2649] == 2649 && 
b[2650] == 2650 && 
b[2651] == 2651 && 
b[2652] == 2652 && 
b[2653] == 2653 && 
b[2654] == 2654 && 
b[2655] == 2655 && 
b[2656] == 2656 && 
b[2657] == 2657 && 
b[2658] == 2658 && 
b[2659] == 2659 && 
b[2660] == 2660 && 
b[2661] == 2661 && 
b[2662] == 2662 && 
b[2663] == 2663 && 
b[2664] == 2664 && 
b[2665] == 2665 && 
b[2666] == 2666 && 
b[2667] == 2667 && 
b[2668] == 2668 && 
b[2669] == 2669 && 
b[2670] == 2670 && 
b[2671] == 2671 && 
b[2672] == 2672 && 
b[2673] == 2673 && 
b[2674] == 2674 && 
b[2675] == 2675 && 
b[2676] == 2676 && 
b[2677] == 2677 && 
b[2678] == 2678 && 
b[2679] == 2679 && 
b[2680] == 2680 && 
b[2681] == 2681 && 
b[2682] == 2682 && 
b[2683] == 2683 && 
b[2684] == 2684 && 
b[2685] == 2685 && 
b[2686] == 2686 && 
b[2687] == 2687 && 
b[2688] == 2688 && 
b[2689] == 2689 && 
b[2690] == 2690 && 
b[2691] == 2691 && 
b[2692] == 2692 && 
b[2693] == 2693 && 
b[2694] == 2694 && 
b[2695] == 2695 && 
b[2696] == 2696 && 
b[2697] == 2697 && 
b[2698] == 2698 && 
b[2699] == 2699 && 
b[2700] == 2700 && 
b[2701] == 2701 && 
b[2702] == 2702 && 
b[2703] == 2703 && 
b[2704] == 2704 && 
b[2705] == 2705 && 
b[2706] == 2706 && 
b[2707] == 2707 && 
b[2708] == 2708 && 
b[2709] == 2709 && 
b[2710] == 2710 && 
b[2711] == 2711 && 
b[2712] == 2712 && 
b[2713] == 2713 && 
b[2714] == 2714 && 
b[2715] == 2715 && 
b[2716] == 2716 && 
b[2717] == 2717 && 
b[2718] == 2718 && 
b[2719] == 2719 && 
b[2720] == 2720 && 
b[2721] == 2721 && 
b[2722] == 2722 && 
b[2723] == 2723 && 
b[2724] == 2724 && 
b[2725] == 2725 && 
b[2726] == 2726 && 
b[2727] == 2727 && 
b[2728] == 2728 && 
b[2729] == 2729 && 
b[2730] == 2730 && 
b[2731] == 2731 && 
b[2732] == 2732 && 
b[2733] == 2733 && 
b[2734] == 2734 && 
b[2735] == 2735 && 
b[2736] == 2736 && 
b[2737] == 2737 && 
b[2738] == 2738 && 
b[2739] == 2739 && 
b[2740] == 2740 && 
b[2741] == 2741 && 
b[2742] == 2742 && 
b[2743] == 2743 && 
b[2744] == 2744 && 
b[2745] == 2745 && 
b[2746] == 2746 && 
b[2747] == 2747 && 
b[2748] == 2748 && 
b[2749] == 2749 && 
b[2750] == 2750 && 
b[2751] == 2751 && 
b[2752] == 2752 && 
b[2753] == 2753 && 
b[2754] == 2754 && 
b[2755] == 2755 && 
b[2756] == 2756 && 
b[2757] == 2757 && 
b[2758] == 2758 && 
b[2759] == 2759 && 
b[2760] == 2760 && 
b[2761] == 2761 && 
b[2762] == 2762 && 
b[2763] == 2763 && 
b[2764] == 2764 && 
b[2765] == 2765 && 
b[2766] == 2766 && 
b[2767] == 2767 && 
b[2768] == 2768 && 
b[2769] == 2769 && 
b[2770] == 2770 && 
b[2771] == 2771 && 
b[2772] == 2772 && 
b[2773] == 2773 && 
b[2774] == 2774 && 
b[2775] == 2775 && 
b[2776] == 2776 && 
b[2777] == 2777 && 
b[2778] == 2778 && 
b[2779] == 2779 && 
b[2780] == 2780 && 
b[2781] == 2781 && 
b[2782] == 2782 && 
b[2783] == 2783 && 
b[2784] == 2784 && 
b[2785] == 2785 && 
b[2786] == 2786 && 
b[2787] == 2787 && 
b[2788] == 2788 && 
b[2789] == 2789 && 
b[2790] == 2790 && 
b[2791] == 2791 && 
b[2792] == 2792 && 
b[2793] == 2793 && 
b[2794] == 2794 && 
b[2795] == 2795 && 
b[2796] == 2796 && 
b[2797] == 2797 && 
b[2798] == 2798 && 
b[2799] == 2799 && 
b[2800] == 2800 && 
b[2801] == 2801 && 
b[2802] == 2802 && 
b[2803] == 2803 && 
b[2804] == 2804 && 
b[2805] == 2805 && 
b[2806] == 2806 && 
b[2807] == 2807 && 
b[2808] == 2808 && 
b[2809] == 2809 && 
b[2810] == 2810 && 
b[2811] == 2811 && 
b[2812] == 2812 && 
b[2813] == 2813 && 
b[2814] == 2814 && 
b[2815] == 2815 && 
b[2816] == 2816 && 
b[2817] == 2817 && 
b[2818] == 2818 && 
b[2819] == 2819 && 
b[2820] == 2820 && 
b[2821] == 2821 && 
b[2822] == 2822 && 
b[2823] == 2823 && 
b[2824] == 2824 && 
b[2825] == 2825 && 
b[2826] == 2826 && 
b[2827] == 2827 && 
b[2828] == 2828 && 
b[2829] == 2829 && 
b[2830] == 2830 && 
b[2831] == 2831 && 
b[2832] == 2832 && 
b[2833] == 2833 && 
b[2834] == 2834 && 
b[2835] == 2835 && 
b[2836] == 2836 && 
b[2837] == 2837 && 
b[2838] == 2838 && 
b[2839] == 2839 && 
b[2840] == 2840 && 
b[2841] == 2841 && 
b[2842] == 2842 && 
b[2843] == 2843 && 
b[2844] == 2844 && 
b[2845] == 2845 && 
b[2846] == 2846 && 
b[2847] == 2847 && 
b[2848] == 2848 && 
b[2849] == 2849 && 
b[2850] == 2850 && 
b[2851] == 2851 && 
b[2852] == 2852 && 
b[2853] == 2853 && 
b[2854] == 2854 && 
b[2855] == 2855 && 
b[2856] == 2856 && 
b[2857] == 2857 && 
b[2858] == 2858 && 
b[2859] == 2859 && 
b[2860] == 2860 && 
b[2861] == 2861 && 
b[2862] == 2862 && 
b[2863] == 2863 && 
b[2864] == 2864 && 
b[2865] == 2865 && 
b[2866] == 2866 && 
b[2867] == 2867 && 
b[2868] == 2868 && 
b[2869] == 2869 && 
b[2870] == 2870 && 
b[2871] == 2871 && 
b[2872] == 2872 && 
b[2873] == 2873 && 
b[2874] == 2874 && 
b[2875] == 2875 && 
b[2876] == 2876 && 
b[2877] == 2877 && 
b[2878] == 2878 && 
b[2879] == 2879 && 
b[2880] == 2880 && 
b[2881] == 2881 && 
b[2882] == 2882 && 
b[2883] == 2883 && 
b[2884] == 2884 && 
b[2885] == 2885 && 
b[2886] == 2886 && 
b[2887] == 2887 && 
b[2888] == 2888 && 
b[2889] == 2889 && 
b[2890] == 2890 && 
b[2891] == 2891 && 
b[2892] == 2892 && 
b[2893] == 2893 && 
b[2894] == 2894 && 
b[2895] == 2895 && 
b[2896] == 2896 && 
b[2897] == 2897 && 
b[2898] == 2898 && 
b[2899] == 2899 && 
b[2900] == 2900 && 
b[2901] == 2901 && 
b[2902] == 2902 && 
b[2903] == 2903 && 
b[2904] == 2904 && 
b[2905] == 2905 && 
b[2906] == 2906 && 
b[2907] == 2907 && 
b[2908] == 2908 && 
b[2909] == 2909 && 
b[2910] == 2910 && 
b[2911] == 2911 && 
b[2912] == 2912 && 
b[2913] == 2913 && 
b[2914] == 2914 && 
b[2915] == 2915 && 
b[2916] == 2916 && 
b[2917] == 2917 && 
b[2918] == 2918 && 
b[2919] == 2919 && 
b[2920] == 2920 && 
b[2921] == 2921 && 
b[2922] == 2922 && 
b[2923] == 2923 && 
b[2924] == 2924 && 
b[2925] == 2925 && 
b[2926] == 2926 && 
b[2927] == 2927 && 
b[2928] == 2928 && 
b[2929] == 2929 && 
b[2930] == 2930 && 
b[2931] == 2931 && 
b[2932] == 2932 && 
b[2933] == 2933 && 
b[2934] == 2934 && 
b[2935] == 2935 && 
b[2936] == 2936 && 
b[2937] == 2937 && 
b[2938] == 2938 && 
b[2939] == 2939 && 
b[2940] == 2940 && 
b[2941] == 2941 && 
b[2942] == 2942 && 
b[2943] == 2943 && 
b[2944] == 2944 && 
b[2945] == 2945 && 
b[2946] == 2946 && 
b[2947] == 2947 && 
b[2948] == 2948 && 
b[2949] == 2949 && 
b[2950] == 2950 && 
b[2951] == 2951 && 
b[2952] == 2952 && 
b[2953] == 2953 && 
b[2954] == 2954 && 
b[2955] == 2955 && 
b[2956] == 2956 && 
b[2957] == 2957 && 
b[2958] == 2958 && 
b[2959] == 2959 && 
b[2960] == 2960 && 
b[2961] == 2961 && 
b[2962] == 2962 && 
b[2963] == 2963 && 
b[2964] == 2964 && 
b[2965] == 2965 && 
b[2966] == 2966 && 
b[2967] == 2967 && 
b[2968] == 2968 && 
b[2969] == 2969 && 
b[2970] == 2970 && 
b[2971] == 2971 && 
b[2972] == 2972 && 
b[2973] == 2973 && 
b[2974] == 2974 && 
b[2975] == 2975 && 
b[2976] == 2976 && 
b[2977] == 2977 && 
b[2978] == 2978 && 
b[2979] == 2979 && 
b[2980] == 2980 && 
b[2981] == 2981 && 
b[2982] == 2982 && 
b[2983] == 2983 && 
b[2984] == 2984 && 
b[2985] == 2985 && 
b[2986] == 2986 && 
b[2987] == 2987 && 
b[2988] == 2988 && 
b[2989] == 2989 && 
b[2990] == 2990 && 
b[2991] == 2991 && 
b[2992] == 2992 && 
b[2993] == 2993 && 
b[2994] == 2994 && 
b[2995] == 2995 && 
b[2996] == 2996 && 
b[2997] == 2997 && 
b[2998] == 2998 && 
b[2999] == 2999 && 
b[3000] == 3000 && 
b[3001] == 3001 && 
b[3002] == 3002 && 
b[3003] == 3003 && 
b[3004] == 3004 && 
b[3005] == 3005 && 
b[3006] == 3006 && 
b[3007] == 3007 && 
b[3008] == 3008 && 
b[3009] == 3009 && 
b[3010] == 3010 && 
b[3011] == 3011 && 
b[3012] == 3012 && 
b[3013] == 3013 && 
b[3014] == 3014 && 
b[3015] == 3015 && 
b[3016] == 3016 && 
b[3017] == 3017 && 
b[3018] == 3018 && 
b[3019] == 3019 && 
b[3020] == 3020 && 
b[3021] == 3021 && 
b[3022] == 3022 && 
b[3023] == 3023 && 
b[3024] == 3024 && 
b[3025] == 3025 && 
b[3026] == 3026 && 
b[3027] == 3027 && 
b[3028] == 3028 && 
b[3029] == 3029 && 
b[3030] == 3030 && 
b[3031] == 3031 && 
b[3032] == 3032 && 
b[3033] == 3033 && 
b[3034] == 3034 && 
b[3035] == 3035 && 
b[3036] == 3036 && 
b[3037] == 3037 && 
b[3038] == 3038 && 
b[3039] == 3039 && 
b[3040] == 3040 && 
b[3041] == 3041 && 
b[3042] == 3042 && 
b[3043] == 3043 && 
b[3044] == 3044 && 
b[3045] == 3045 && 
b[3046] == 3046 && 
b[3047] == 3047 && 
b[3048] == 3048 && 
b[3049] == 3049 && 
b[3050] == 3050 && 
b[3051] == 3051 && 
b[3052] == 3052 && 
b[3053] == 3053 && 
b[3054] == 3054 && 
b[3055] == 3055 && 
b[3056] == 3056 && 
b[3057] == 3057 && 
b[3058] == 3058 && 
b[3059] == 3059 && 
b[3060] == 3060 && 
b[3061] == 3061 && 
b[3062] == 3062 && 
b[3063] == 3063 && 
b[3064] == 3064 && 
b[3065] == 3065 && 
b[3066] == 3066 && 
b[3067] == 3067 && 
b[3068] == 3068 && 
b[3069] == 3069 && 
b[3070] == 3070 && 
b[3071] == 3071 && 
b[3072] == 3072 && 
b[3073] == 3073 && 
b[3074] == 3074 && 
b[3075] == 3075 && 
b[3076] == 3076 && 
b[3077] == 3077 && 
b[3078] == 3078 && 
b[3079] == 3079 && 
b[3080] == 3080 && 
b[3081] == 3081 && 
b[3082] == 3082 && 
b[3083] == 3083 && 
b[3084] == 3084 && 
b[3085] == 3085 && 
b[3086] == 3086 && 
b[3087] == 3087 && 
b[3088] == 3088 && 
b[3089] == 3089 && 
b[3090] == 3090 && 
b[3091] == 3091 && 
b[3092] == 3092 && 
b[3093] == 3093 && 
b[3094] == 3094 && 
b[3095] == 3095 && 
b[3096] == 3096 && 
b[3097] == 3097 && 
b[3098] == 3098 && 
b[3099] == 3099 && 
b[3100] == 3100 && 
b[3101] == 3101 && 
b[3102] == 3102 && 
b[3103] == 3103 && 
b[3104] == 3104 && 
b[3105] == 3105 && 
b[3106] == 3106 && 
b[3107] == 3107 && 
b[3108] == 3108 && 
b[3109] == 3109 && 
b[3110] == 3110 && 
b[3111] == 3111 && 
b[3112] == 3112 && 
b[3113] == 3113 && 
b[3114] == 3114 && 
b[3115] == 3115 && 
b[3116] == 3116 && 
b[3117] == 3117 && 
b[3118] == 3118 && 
b[3119] == 3119 && 
b[3120] == 3120 && 
b[3121] == 3121 && 
b[3122] == 3122 && 
b[3123] == 3123 && 
b[3124] == 3124 && 
b[3125] == 3125 && 
b[3126] == 3126 && 
b[3127] == 3127 && 
b[3128] == 3128 && 
b[3129] == 3129 && 
b[3130] == 3130 && 
b[3131] == 3131 && 
b[3132] == 3132 && 
b[3133] == 3133 && 
b[3134] == 3134 && 
b[3135] == 3135 && 
b[3136] == 3136 && 
b[3137] == 3137 && 
b[3138] == 3138 && 
b[3139] == 3139 && 
b[3140] == 3140 && 
b[3141] == 3141 && 
b[3142] == 3142 && 
b[3143] == 3143 && 
b[3144] == 3144 && 
b[3145] == 3145 && 
b[3146] == 3146 && 
b[3147] == 3147 && 
b[3148] == 3148 && 
b[3149] == 3149 && 
b[3150] == 3150 && 
b[3151] == 3151 && 
b[3152] == 3152 && 
b[3153] == 3153 && 
b[3154] == 3154 && 
b[3155] == 3155 && 
b[3156] == 3156 && 
b[3157] == 3157 && 
b[3158] == 3158 && 
b[3159] == 3159 && 
b[3160] == 3160 && 
b[3161] == 3161 && 
b[3162] == 3162 && 
b[3163] == 3163 && 
b[3164] == 3164 && 
b[3165] == 3165 && 
b[3166] == 3166 && 
b[3167] == 3167 && 
b[3168] == 3168 && 
b[3169] == 3169 && 
b[3170] == 3170 && 
b[3171] == 3171 && 
b[3172] == 3172 && 
b[3173] == 3173 && 
b[3174] == 3174 && 
b[3175] == 3175 && 
b[3176] == 3176 && 
b[3177] == 3177 && 
b[3178] == 3178 && 
b[3179] == 3179 && 
b[3180] == 3180 && 
b[3181] == 3181 && 
b[3182] == 3182 && 
b[3183] == 3183 && 
b[3184] == 3184 && 
b[3185] == 3185 && 
b[3186] == 3186 && 
b[3187] == 3187 && 
b[3188] == 3188 && 
b[3189] == 3189 && 
b[3190] == 3190 && 
b[3191] == 3191 && 
b[3192] == 3192 && 
b[3193] == 3193 && 
b[3194] == 3194 && 
b[3195] == 3195 && 
b[3196] == 3196 && 
b[3197] == 3197 && 
b[3198] == 3198 && 
b[3199] == 3199 && 
b[3200] == 3200 && 
b[3201] == 3201 && 
b[3202] == 3202 && 
b[3203] == 3203 && 
b[3204] == 3204 && 
b[3205] == 3205 && 
b[3206] == 3206 && 
b[3207] == 3207 && 
b[3208] == 3208 && 
b[3209] == 3209 && 
b[3210] == 3210 && 
b[3211] == 3211 && 
b[3212] == 3212 && 
b[3213] == 3213 && 
b[3214] == 3214 && 
b[3215] == 3215 && 
b[3216] == 3216 && 
b[3217] == 3217 && 
b[3218] == 3218 && 
b[3219] == 3219 && 
b[3220] == 3220 && 
b[3221] == 3221 && 
b[3222] == 3222 && 
b[3223] == 3223 && 
b[3224] == 3224 && 
b[3225] == 3225 && 
b[3226] == 3226 && 
b[3227] == 3227 && 
b[3228] == 3228 && 
b[3229] == 3229 && 
b[3230] == 3230 && 
b[3231] == 3231 && 
b[3232] == 3232 && 
b[3233] == 3233 && 
b[3234] == 3234 && 
b[3235] == 3235 && 
b[3236] == 3236 && 
b[3237] == 3237 && 
b[3238] == 3238 && 
b[3239] == 3239 && 
b[3240] == 3240 && 
b[3241] == 3241 && 
b[3242] == 3242 && 
b[3243] == 3243 && 
b[3244] == 3244 && 
b[3245] == 3245 && 
b[3246] == 3246 && 
b[3247] == 3247 && 
b[3248] == 3248 && 
b[3249] == 3249 && 
b[3250] == 3250 && 
b[3251] == 3251 && 
b[3252] == 3252 && 
b[3253] == 3253 && 
b[3254] == 3254 && 
b[3255] == 3255 && 
b[3256] == 3256 && 
b[3257] == 3257 && 
b[3258] == 3258 && 
b[3259] == 3259 && 
b[3260] == 3260 && 
b[3261] == 3261 && 
b[3262] == 3262 && 
b[3263] == 3263 && 
b[3264] == 3264 && 
b[3265] == 3265 && 
b[3266] == 3266 && 
b[3267] == 3267 && 
b[3268] == 3268 && 
b[3269] == 3269 && 
b[3270] == 3270 && 
b[3271] == 3271 && 
b[3272] == 3272 && 
b[3273] == 3273 && 
b[3274] == 3274 && 
b[3275] == 3275 && 
b[3276] == 3276 && 
b[3277] == 3277 && 
b[3278] == 3278 && 
b[3279] == 3279 && 
b[3280] == 3280 && 
b[3281] == 3281 && 
b[3282] == 3282 && 
b[3283] == 3283 && 
b[3284] == 3284 && 
b[3285] == 3285 && 
b[3286] == 3286 && 
b[3287] == 3287 && 
b[3288] == 3288 && 
b[3289] == 3289 && 
b[3290] == 3290 && 
b[3291] == 3291 && 
b[3292] == 3292 && 
b[3293] == 3293 && 
b[3294] == 3294 && 
b[3295] == 3295 && 
b[3296] == 3296 && 
b[3297] == 3297 && 
b[3298] == 3298 && 
b[3299] == 3299 && 
b[3300] == 3300 && 
b[3301] == 3301 && 
b[3302] == 3302 && 
b[3303] == 3303 && 
b[3304] == 3304 && 
b[3305] == 3305 && 
b[3306] == 3306 && 
b[3307] == 3307 && 
b[3308] == 3308 && 
b[3309] == 3309 && 
b[3310] == 3310 && 
b[3311] == 3311 && 
b[3312] == 3312 && 
b[3313] == 3313 && 
b[3314] == 3314 && 
b[3315] == 3315 && 
b[3316] == 3316 && 
b[3317] == 3317 && 
b[3318] == 3318 && 
b[3319] == 3319 && 
b[3320] == 3320 && 
b[3321] == 3321 && 
b[3322] == 3322 && 
b[3323] == 3323 && 
b[3324] == 3324 && 
b[3325] == 3325 && 
b[3326] == 3326 && 
b[3327] == 3327 && 
b[3328] == 3328 && 
b[3329] == 3329 && 
b[3330] == 3330 && 
b[3331] == 3331 && 
b[3332] == 3332 && 
b[3333] == 3333 && 
b[3334] == 3334 && 
b[3335] == 3335 && 
b[3336] == 3336 && 
b[3337] == 3337 && 
b[3338] == 3338 && 
b[3339] == 3339 && 
b[3340] == 3340 && 
b[3341] == 3341 && 
b[3342] == 3342 && 
b[3343] == 3343 && 
b[3344] == 3344 && 
b[3345] == 3345 && 
b[3346] == 3346 && 
b[3347] == 3347 && 
b[3348] == 3348 && 
b[3349] == 3349 && 
b[3350] == 3350 && 
b[3351] == 3351 && 
b[3352] == 3352 && 
b[3353] == 3353 && 
b[3354] == 3354 && 
b[3355] == 3355 && 
b[3356] == 3356 && 
b[3357] == 3357 && 
b[3358] == 3358 && 
b[3359] == 3359 && 
b[3360] == 3360 && 
b[3361] == 3361 && 
b[3362] == 3362 && 
b[3363] == 3363 && 
b[3364] == 3364 && 
b[3365] == 3365 && 
b[3366] == 3366 && 
b[3367] == 3367 && 
b[3368] == 3368 && 
b[3369] == 3369 && 
b[3370] == 3370 && 
b[3371] == 3371 && 
b[3372] == 3372 && 
b[3373] == 3373 && 
b[3374] == 3374 && 
b[3375] == 3375 && 
b[3376] == 3376 && 
b[3377] == 3377 && 
b[3378] == 3378 && 
b[3379] == 3379 && 
b[3380] == 3380 && 
b[3381] == 3381 && 
b[3382] == 3382 && 
b[3383] == 3383 && 
b[3384] == 3384 && 
b[3385] == 3385 && 
b[3386] == 3386 && 
b[3387] == 3387 && 
b[3388] == 3388 && 
b[3389] == 3389 && 
b[3390] == 3390 && 
b[3391] == 3391 && 
b[3392] == 3392 && 
b[3393] == 3393 && 
b[3394] == 3394 && 
b[3395] == 3395 && 
b[3396] == 3396 && 
b[3397] == 3397 && 
b[3398] == 3398 && 
b[3399] == 3399 && 
b[3400] == 3400 && 
b[3401] == 3401 && 
b[3402] == 3402 && 
b[3403] == 3403 && 
b[3404] == 3404 && 
b[3405] == 3405 && 
b[3406] == 3406 && 
b[3407] == 3407 && 
b[3408] == 3408 && 
b[3409] == 3409 && 
b[3410] == 3410 && 
b[3411] == 3411 && 
b[3412] == 3412 && 
b[3413] == 3413 && 
b[3414] == 3414 && 
b[3415] == 3415 && 
b[3416] == 3416 && 
b[3417] == 3417 && 
b[3418] == 3418 && 
b[3419] == 3419 && 
b[3420] == 3420 && 
b[3421] == 3421 && 
b[3422] == 3422 && 
b[3423] == 3423 && 
b[3424] == 3424 && 
b[3425] == 3425 && 
b[3426] == 3426 && 
b[3427] == 3427 && 
b[3428] == 3428 && 
b[3429] == 3429 && 
b[3430] == 3430 && 
b[3431] == 3431 && 
b[3432] == 3432 && 
b[3433] == 3433 && 
b[3434] == 3434 && 
b[3435] == 3435 && 
b[3436] == 3436 && 
b[3437] == 3437 && 
b[3438] == 3438 && 
b[3439] == 3439 && 
b[3440] == 3440 && 
b[3441] == 3441 && 
b[3442] == 3442 && 
b[3443] == 3443 && 
b[3444] == 3444 && 
b[3445] == 3445 && 
b[3446] == 3446 && 
b[3447] == 3447 && 
b[3448] == 3448 && 
b[3449] == 3449 && 
b[3450] == 3450 && 
b[3451] == 3451 && 
b[3452] == 3452 && 
b[3453] == 3453 && 
b[3454] == 3454 && 
b[3455] == 3455 && 
b[3456] == 3456 && 
b[3457] == 3457 && 
b[3458] == 3458 && 
b[3459] == 3459 && 
b[3460] == 3460 && 
b[3461] == 3461 && 
b[3462] == 3462 && 
b[3463] == 3463 && 
b[3464] == 3464 && 
b[3465] == 3465 && 
b[3466] == 3466 && 
b[3467] == 3467 && 
b[3468] == 3468 && 
b[3469] == 3469 && 
b[3470] == 3470 && 
b[3471] == 3471 && 
b[3472] == 3472 && 
b[3473] == 3473 && 
b[3474] == 3474 && 
b[3475] == 3475 && 
b[3476] == 3476 && 
b[3477] == 3477 && 
b[3478] == 3478 && 
b[3479] == 3479 && 
b[3480] == 3480 && 
b[3481] == 3481 && 
b[3482] == 3482 && 
b[3483] == 3483 && 
b[3484] == 3484 && 
b[3485] == 3485 && 
b[3486] == 3486 && 
b[3487] == 3487 && 
b[3488] == 3488 && 
b[3489] == 3489 && 
b[3490] == 3490 && 
b[3491] == 3491 && 
b[3492] == 3492 && 
b[3493] == 3493 && 
b[3494] == 3494 && 
b[3495] == 3495 && 
b[3496] == 3496 && 
b[3497] == 3497 && 
b[3498] == 3498 && 
b[3499] == 3499 && 
b[3500] == 3500 && 
b[3501] == 3501 && 
b[3502] == 3502 && 
b[3503] == 3503 && 
b[3504] == 3504 && 
b[3505] == 3505 && 
b[3506] == 3506 && 
b[3507] == 3507 && 
b[3508] == 3508 && 
b[3509] == 3509 && 
b[3510] == 3510 && 
b[3511] == 3511 && 
b[3512] == 3512 && 
b[3513] == 3513 && 
b[3514] == 3514 && 
b[3515] == 3515 && 
b[3516] == 3516 && 
b[3517] == 3517 && 
b[3518] == 3518 && 
b[3519] == 3519 && 
b[3520] == 3520 && 
b[3521] == 3521 && 
b[3522] == 3522 && 
b[3523] == 3523 && 
b[3524] == 3524 && 
b[3525] == 3525 && 
b[3526] == 3526 && 
b[3527] == 3527 && 
b[3528] == 3528 && 
b[3529] == 3529 && 
b[3530] == 3530 && 
b[3531] == 3531 && 
b[3532] == 3532 && 
b[3533] == 3533 && 
b[3534] == 3534 && 
b[3535] == 3535 && 
b[3536] == 3536 && 
b[3537] == 3537 && 
b[3538] == 3538 && 
b[3539] == 3539 && 
b[3540] == 3540 && 
b[3541] == 3541 && 
b[3542] == 3542 && 
b[3543] == 3543 && 
b[3544] == 3544 && 
b[3545] == 3545 && 
b[3546] == 3546 && 
b[3547] == 3547 && 
b[3548] == 3548 && 
b[3549] == 3549 && 
b[3550] == 3550 && 
b[3551] == 3551 && 
b[3552] == 3552 && 
b[3553] == 3553 && 
b[3554] == 3554 && 
b[3555] == 3555 && 
b[3556] == 3556 && 
b[3557] == 3557 && 
b[3558] == 3558 && 
b[3559] == 3559 && 
b[3560] == 3560 && 
b[3561] == 3561 && 
b[3562] == 3562 && 
b[3563] == 3563 && 
b[3564] == 3564 && 
b[3565] == 3565 && 
b[3566] == 3566 && 
b[3567] == 3567 && 
b[3568] == 3568 && 
b[3569] == 3569 && 
b[3570] == 3570 && 
b[3571] == 3571 && 
b[3572] == 3572 && 
b[3573] == 3573 && 
b[3574] == 3574 && 
b[3575] == 3575 && 
b[3576] == 3576 && 
b[3577] == 3577 && 
b[3578] == 3578 && 
b[3579] == 3579 && 
b[3580] == 3580 && 
b[3581] == 3581 && 
b[3582] == 3582 && 
b[3583] == 3583 && 
b[3584] == 3584 && 
b[3585] == 3585 && 
b[3586] == 3586 && 
b[3587] == 3587 && 
b[3588] == 3588 && 
b[3589] == 3589 && 
b[3590] == 3590 && 
b[3591] == 3591 && 
b[3592] == 3592 && 
b[3593] == 3593 && 
b[3594] == 3594 && 
b[3595] == 3595 && 
b[3596] == 3596 && 
b[3597] == 3597 && 
b[3598] == 3598 && 
b[3599] == 3599 && 
b[3600] == 3600 && 
b[3601] == 3601 && 
b[3602] == 3602 && 
b[3603] == 3603 && 
b[3604] == 3604 && 
b[3605] == 3605 && 
b[3606] == 3606 && 
b[3607] == 3607 && 
b[3608] == 3608 && 
b[3609] == 3609 && 
b[3610] == 3610 && 
b[3611] == 3611 && 
b[3612] == 3612 && 
b[3613] == 3613 && 
b[3614] == 3614 && 
b[3615] == 3615 && 
b[3616] == 3616 && 
b[3617] == 3617 && 
b[3618] == 3618 && 
b[3619] == 3619 && 
b[3620] == 3620 && 
b[3621] == 3621 && 
b[3622] == 3622 && 
b[3623] == 3623 && 
b[3624] == 3624 && 
b[3625] == 3625 && 
b[3626] == 3626 && 
b[3627] == 3627 && 
b[3628] == 3628 && 
b[3629] == 3629 && 
b[3630] == 3630 && 
b[3631] == 3631 && 
b[3632] == 3632 && 
b[3633] == 3633 && 
b[3634] == 3634 && 
b[3635] == 3635 && 
b[3636] == 3636 && 
b[3637] == 3637 && 
b[3638] == 3638 && 
b[3639] == 3639 && 
b[3640] == 3640 && 
b[3641] == 3641 && 
b[3642] == 3642 && 
b[3643] == 3643 && 
b[3644] == 3644 && 
b[3645] == 3645 && 
b[3646] == 3646 && 
b[3647] == 3647 && 
b[3648] == 3648 && 
b[3649] == 3649 && 
b[3650] == 3650 && 
b[3651] == 3651 && 
b[3652] == 3652 && 
b[3653] == 3653 && 
b[3654] == 3654 && 
b[3655] == 3655 && 
b[3656] == 3656 && 
b[3657] == 3657 && 
b[3658] == 3658 && 
b[3659] == 3659 && 
b[3660] == 3660 && 
b[3661] == 3661 && 
b[3662] == 3662 && 
b[3663] == 3663 && 
b[3664] == 3664 && 
b[3665] == 3665 && 
b[3666] == 3666 && 
b[3667] == 3667 && 
b[3668] == 3668 && 
b[3669] == 3669 && 
b[3670] == 3670 && 
b[3671] == 3671 && 
b[3672] == 3672 && 
b[3673] == 3673 && 
b[3674] == 3674 && 
b[3675] == 3675 && 
b[3676] == 3676 && 
b[3677] == 3677 && 
b[3678] == 3678 && 
b[3679] == 3679 && 
b[3680] == 3680 && 
b[3681] == 3681 && 
b[3682] == 3682 && 
b[3683] == 3683 && 
b[3684] == 3684 && 
b[3685] == 3685 && 
b[3686] == 3686 && 
b[3687] == 3687 && 
b[3688] == 3688 && 
b[3689] == 3689 && 
b[3690] == 3690 && 
b[3691] == 3691 && 
b[3692] == 3692 && 
b[3693] == 3693 && 
b[3694] == 3694 && 
b[3695] == 3695 && 
b[3696] == 3696 && 
b[3697] == 3697 && 
b[3698] == 3698 && 
b[3699] == 3699 && 
b[3700] == 3700 && 
b[3701] == 3701 && 
b[3702] == 3702 && 
b[3703] == 3703 && 
b[3704] == 3704 && 
b[3705] == 3705 && 
b[3706] == 3706 && 
b[3707] == 3707 && 
b[3708] == 3708 && 
b[3709] == 3709 && 
b[3710] == 3710 && 
b[3711] == 3711 && 
b[3712] == 3712 && 
b[3713] == 3713 && 
b[3714] == 3714 && 
b[3715] == 3715 && 
b[3716] == 3716 && 
b[3717] == 3717 && 
b[3718] == 3718 && 
b[3719] == 3719 && 
b[3720] == 3720 && 
b[3721] == 3721 && 
b[3722] == 3722 && 
b[3723] == 3723 && 
b[3724] == 3724 && 
b[3725] == 3725 && 
b[3726] == 3726 && 
b[3727] == 3727 && 
b[3728] == 3728 && 
b[3729] == 3729 && 
b[3730] == 3730 && 
b[3731] == 3731 && 
b[3732] == 3732 && 
b[3733] == 3733 && 
b[3734] == 3734 && 
b[3735] == 3735 && 
b[3736] == 3736 && 
b[3737] == 3737 && 
b[3738] == 3738 && 
b[3739] == 3739 && 
b[3740] == 3740 && 
b[3741] == 3741 && 
b[3742] == 3742 && 
b[3743] == 3743 && 
b[3744] == 3744 && 
b[3745] == 3745 && 
b[3746] == 3746 && 
b[3747] == 3747 && 
b[3748] == 3748 && 
b[3749] == 3749 && 
b[3750] == 3750 && 
b[3751] == 3751 && 
b[3752] == 3752 && 
b[3753] == 3753 && 
b[3754] == 3754 && 
b[3755] == 3755 && 
b[3756] == 3756 && 
b[3757] == 3757 && 
b[3758] == 3758 && 
b[3759] == 3759 && 
b[3760] == 3760 && 
b[3761] == 3761 && 
b[3762] == 3762 && 
b[3763] == 3763 && 
b[3764] == 3764 && 
b[3765] == 3765 && 
b[3766] == 3766 && 
b[3767] == 3767 && 
b[3768] == 3768 && 
b[3769] == 3769 && 
b[3770] == 3770 && 
b[3771] == 3771 && 
b[3772] == 3772 && 
b[3773] == 3773 && 
b[3774] == 3774 && 
b[3775] == 3775 && 
b[3776] == 3776 && 
b[3777] == 3777 && 
b[3778] == 3778 && 
b[3779] == 3779 && 
b[3780] == 3780 && 
b[3781] == 3781 && 
b[3782] == 3782 && 
b[3783] == 3783 && 
b[3784] == 3784 && 
b[3785] == 3785 && 
b[3786] == 3786 && 
b[3787] == 3787 && 
b[3788] == 3788 && 
b[3789] == 3789 && 
b[3790] == 3790 && 
b[3791] == 3791 && 
b[3792] == 3792 && 
b[3793] == 3793 && 
b[3794] == 3794 && 
b[3795] == 3795 && 
b[3796] == 3796 && 
b[3797] == 3797 && 
b[3798] == 3798 && 
b[3799] == 3799 && 
b[3800] == 3800 && 
b[3801] == 3801 && 
b[3802] == 3802 && 
b[3803] == 3803 && 
b[3804] == 3804 && 
b[3805] == 3805 && 
b[3806] == 3806 && 
b[3807] == 3807 && 
b[3808] == 3808 && 
b[3809] == 3809 && 
b[3810] == 3810 && 
b[3811] == 3811 && 
b[3812] == 3812 && 
b[3813] == 3813 && 
b[3814] == 3814 && 
b[3815] == 3815 && 
b[3816] == 3816 && 
b[3817] == 3817 && 
b[3818] == 3818 && 
b[3819] == 3819 && 
b[3820] == 3820 && 
b[3821] == 3821 && 
b[3822] == 3822 && 
b[3823] == 3823 && 
b[3824] == 3824 && 
b[3825] == 3825 && 
b[3826] == 3826 && 
b[3827] == 3827 && 
b[3828] == 3828 && 
b[3829] == 3829 && 
b[3830] == 3830 && 
b[3831] == 3831 && 
b[3832] == 3832 && 
b[3833] == 3833 && 
b[3834] == 3834 && 
b[3835] == 3835 && 
b[3836] == 3836 && 
b[3837] == 3837 && 
b[3838] == 3838 && 
b[3839] == 3839 && 
b[3840] == 3840 && 
b[3841] == 3841 && 
b[3842] == 3842 && 
b[3843] == 3843 && 
b[3844] == 3844 && 
b[3845] == 3845 && 
b[3846] == 3846 && 
b[3847] == 3847 && 
b[3848] == 3848 && 
b[3849] == 3849 && 
b[3850] == 3850 && 
b[3851] == 3851 && 
b[3852] == 3852 && 
b[3853] == 3853 && 
b[3854] == 3854 && 
b[3855] == 3855 && 
b[3856] == 3856 && 
b[3857] == 3857 && 
b[3858] == 3858 && 
b[3859] == 3859 && 
b[3860] == 3860 && 
b[3861] == 3861 && 
b[3862] == 3862 && 
b[3863] == 3863 && 
b[3864] == 3864 && 
b[3865] == 3865 && 
b[3866] == 3866 && 
b[3867] == 3867 && 
b[3868] == 3868 && 
b[3869] == 3869 && 
b[3870] == 3870 && 
b[3871] == 3871 && 
b[3872] == 3872 && 
b[3873] == 3873 && 
b[3874] == 3874 && 
b[3875] == 3875 && 
b[3876] == 3876 && 
b[3877] == 3877 && 
b[3878] == 3878 && 
b[3879] == 3879 && 
b[3880] == 3880 && 
b[3881] == 3881 && 
b[3882] == 3882 && 
b[3883] == 3883 && 
b[3884] == 3884 && 
b[3885] == 3885 && 
b[3886] == 3886 && 
b[3887] == 3887 && 
b[3888] == 3888 && 
b[3889] == 3889 && 
b[3890] == 3890 && 
b[3891] == 3891 && 
b[3892] == 3892 && 
b[3893] == 3893 && 
b[3894] == 3894 && 
b[3895] == 3895 && 
b[3896] == 3896 && 
b[3897] == 3897 && 
b[3898] == 3898 && 
b[3899] == 3899 && 
b[3900] == 3900 && 
b[3901] == 3901 && 
b[3902] == 3902 && 
b[3903] == 3903 && 
b[3904] == 3904 && 
b[3905] == 3905 && 
b[3906] == 3906 && 
b[3907] == 3907 && 
b[3908] == 3908 && 
b[3909] == 3909 && 
b[3910] == 3910 && 
b[3911] == 3911 && 
b[3912] == 3912 && 
b[3913] == 3913 && 
b[3914] == 3914 && 
b[3915] == 3915 && 
b[3916] == 3916 && 
b[3917] == 3917 && 
b[3918] == 3918 && 
b[3919] == 3919 && 
b[3920] == 3920 && 
b[3921] == 3921 && 
b[3922] == 3922 && 
b[3923] == 3923 && 
b[3924] == 3924 && 
b[3925] == 3925 && 
b[3926] == 3926 && 
b[3927] == 3927 && 
b[3928] == 3928 && 
b[3929] == 3929 && 
b[3930] == 3930 && 
b[3931] == 3931 && 
b[3932] == 3932 && 
b[3933] == 3933 && 
b[3934] == 3934 && 
b[3935] == 3935 && 
b[3936] == 3936 && 
b[3937] == 3937 && 
b[3938] == 3938 && 
b[3939] == 3939 && 
b[3940] == 3940 && 
b[3941] == 3941 && 
b[3942] == 3942 && 
b[3943] == 3943 && 
b[3944] == 3944 && 
b[3945] == 3945 && 
b[3946] == 3946 && 
b[3947] == 3947 && 
b[3948] == 3948 && 
b[3949] == 3949 && 
b[3950] == 3950 && 
b[3951] == 3951 && 
b[3952] == 3952 && 
b[3953] == 3953 && 
b[3954] == 3954 && 
b[3955] == 3955 && 
b[3956] == 3956 && 
b[3957] == 3957 && 
b[3958] == 3958 && 
b[3959] == 3959 && 
b[3960] == 3960 && 
b[3961] == 3961 && 
b[3962] == 3962 && 
b[3963] == 3963 && 
b[3964] == 3964 && 
b[3965] == 3965 && 
b[3966] == 3966 && 
b[3967] == 3967 && 
b[3968] == 3968 && 
b[3969] == 3969 && 
b[3970] == 3970 && 
b[3971] == 3971 && 
b[3972] == 3972 && 
b[3973] == 3973 && 
b[3974] == 3974 && 
b[3975] == 3975 && 
b[3976] == 3976 && 
b[3977] == 3977 && 
b[3978] == 3978 && 
b[3979] == 3979 && 
b[3980] == 3980 && 
b[3981] == 3981 && 
b[3982] == 3982 && 
b[3983] == 3983 && 
b[3984] == 3984 && 
b[3985] == 3985 && 
b[3986] == 3986 && 
b[3987] == 3987 && 
b[3988] == 3988 && 
b[3989] == 3989 && 
b[3990] == 3990 && 
b[3991] == 3991 && 
b[3992] == 3992 && 
b[3993] == 3993 && 
b[3994] == 3994 && 
b[3995] == 3995 && 
b[3996] == 3996 && 
b[3997] == 3997 && 
b[3998] == 3998 && 
b[3999] == 3999 && 
b[4000] == 4000 && 
b[4001] == 4001 && 
b[4002] == 4002 && 
b[4003] == 4003 && 
b[4004] == 4004 && 
b[4005] == 4005 && 
b[4006] == 4006 && 
b[4007] == 4007 && 
b[4008] == 4008 && 
b[4009] == 4009 && 
b[4010] == 4010 && 
b[4011] == 4011 && 
b[4012] == 4012 && 
b[4013] == 4013 && 
b[4014] == 4014 && 
b[4015] == 4015 && 
b[4016] == 4016 && 
b[4017] == 4017 && 
b[4018] == 4018 && 
b[4019] == 4019 && 
b[4020] == 4020 && 
b[4021] == 4021 && 
b[4022] == 4022 && 
b[4023] == 4023 && 
b[4024] == 4024 && 
b[4025] == 4025 && 
b[4026] == 4026 && 
b[4027] == 4027 && 
b[4028] == 4028 && 
b[4029] == 4029 && 
b[4030] == 4030 && 
b[4031] == 4031 && 
b[4032] == 4032 && 
b[4033] == 4033 && 
b[4034] == 4034 && 
b[4035] == 4035 && 
b[4036] == 4036 && 
b[4037] == 4037 && 
b[4038] == 4038 && 
b[4039] == 4039 && 
b[4040] == 4040 && 
b[4041] == 4041 && 
b[4042] == 4042 && 
b[4043] == 4043 && 
b[4044] == 4044 && 
b[4045] == 4045 && 
b[4046] == 4046 && 
b[4047] == 4047 && 
b[4048] == 4048 && 
b[4049] == 4049 && 
b[4050] == 4050 && 
b[4051] == 4051 && 
b[4052] == 4052 && 
b[4053] == 4053 && 
b[4054] == 4054 && 
b[4055] == 4055 && 
b[4056] == 4056 && 
b[4057] == 4057 && 
b[4058] == 4058 && 
b[4059] == 4059 && 
b[4060] == 4060 && 
b[4061] == 4061 && 
b[4062] == 4062 && 
b[4063] == 4063 && 
b[4064] == 4064 && 
b[4065] == 4065 && 
b[4066] == 4066 && 
b[4067] == 4067 && 
b[4068] == 4068 && 
b[4069] == 4069 && 
b[4070] == 4070 && 
b[4071] == 4071 && 
b[4072] == 4072 && 
b[4073] == 4073 && 
b[4074] == 4074 && 
b[4075] == 4075 && 
b[4076] == 4076 && 
b[4077] == 4077 && 
b[4078] == 4078 && 
b[4079] == 4079 && 
b[4080] == 4080 && 
b[4081] == 4081 && 
b[4082] == 4082 && 
b[4083] == 4083 && 
b[4084] == 4084 && 
b[4085] == 4085 && 
b[4086] == 4086 && 
b[4087] == 4087 && 
b[4088] == 4088 && 
b[4089] == 4089 && 
b[4090] == 4090 && 
b[4091] == 4091 && 
b[4092] == 4092 && 
b[4093] == 4093 && 
b[4094] == 4094 && 
b[4095] == 4095 && 
b[4096] == 4096 && 
b[4097] == 4097 && 
b[4098] == 4098 && 
b[4099] == 4099 && 
b[4100] == 4100 && 
b[4101] == 4101 && 
b[4102] == 4102 && 
b[4103] == 4103 && 
b[4104] == 4104 && 
b[4105] == 4105 && 
b[4106] == 4106 && 
b[4107] == 4107 && 
b[4108] == 4108 && 
b[4109] == 4109 && 
b[4110] == 4110 && 
b[4111] == 4111 && 
b[4112] == 4112 && 
b[4113] == 4113 && 
b[4114] == 4114 && 
b[4115] == 4115 && 
b[4116] == 4116 && 
b[4117] == 4117 && 
b[4118] == 4118 && 
b[4119] == 4119 && 
b[4120] == 4120 && 
b[4121] == 4121 && 
b[4122] == 4122 && 
b[4123] == 4123 && 
b[4124] == 4124 && 
b[4125] == 4125 && 
b[4126] == 4126 && 
b[4127] == 4127 && 
b[4128] == 4128 && 
b[4129] == 4129 && 
b[4130] == 4130 && 
b[4131] == 4131 && 
b[4132] == 4132 && 
b[4133] == 4133 && 
b[4134] == 4134 && 
b[4135] == 4135 && 
b[4136] == 4136 && 
b[4137] == 4137 && 
b[4138] == 4138 && 
b[4139] == 4139 && 
b[4140] == 4140 && 
b[4141] == 4141 && 
b[4142] == 4142 && 
b[4143] == 4143 && 
b[4144] == 4144 && 
b[4145] == 4145 && 
b[4146] == 4146 && 
b[4147] == 4147 && 
b[4148] == 4148 && 
b[4149] == 4149 && 
b[4150] == 4150 && 
b[4151] == 4151 && 
b[4152] == 4152 && 
b[4153] == 4153 && 
b[4154] == 4154 && 
b[4155] == 4155 && 
b[4156] == 4156 && 
b[4157] == 4157 && 
b[4158] == 4158 && 
b[4159] == 4159 && 
b[4160] == 4160 && 
b[4161] == 4161 && 
b[4162] == 4162 && 
b[4163] == 4163 && 
b[4164] == 4164 && 
b[4165] == 4165 && 
b[4166] == 4166 && 
b[4167] == 4167 && 
b[4168] == 4168 && 
b[4169] == 4169 && 
b[4170] == 4170 && 
b[4171] == 4171 && 
b[4172] == 4172 && 
b[4173] == 4173 && 
b[4174] == 4174 && 
b[4175] == 4175 && 
b[4176] == 4176 && 
b[4177] == 4177 && 
b[4178] == 4178 && 
b[4179] == 4179 && 
b[4180] == 4180 && 
b[4181] == 4181 && 
b[4182] == 4182 && 
b[4183] == 4183 && 
b[4184] == 4184 && 
b[4185] == 4185 && 
b[4186] == 4186 && 
b[4187] == 4187 && 
b[4188] == 4188 && 
b[4189] == 4189 && 
b[4190] == 4190 && 
b[4191] == 4191 && 
b[4192] == 4192 && 
b[4193] == 4193 && 
b[4194] == 4194 && 
b[4195] == 4195 && 
b[4196] == 4196 && 
b[4197] == 4197 && 
b[4198] == 4198 && 
b[4199] == 4199 && 
b[4200] == 4200 && 
b[4201] == 4201 && 
b[4202] == 4202 && 
b[4203] == 4203 && 
b[4204] == 4204 && 
b[4205] == 4205 && 
b[4206] == 4206 && 
b[4207] == 4207 && 
b[4208] == 4208 && 
b[4209] == 4209 && 
b[4210] == 4210 && 
b[4211] == 4211 && 
b[4212] == 4212 && 
b[4213] == 4213 && 
b[4214] == 4214 && 
b[4215] == 4215 && 
b[4216] == 4216 && 
b[4217] == 4217 && 
b[4218] == 4218 && 
b[4219] == 4219 && 
b[4220] == 4220 && 
b[4221] == 4221 && 
b[4222] == 4222 && 
b[4223] == 4223 && 
b[4224] == 4224 && 
b[4225] == 4225 && 
b[4226] == 4226 && 
b[4227] == 4227 && 
b[4228] == 4228 && 
b[4229] == 4229 && 
b[4230] == 4230 && 
b[4231] == 4231 && 
b[4232] == 4232 && 
b[4233] == 4233 && 
b[4234] == 4234 && 
b[4235] == 4235 && 
b[4236] == 4236 && 
b[4237] == 4237 && 
b[4238] == 4238 && 
b[4239] == 4239 && 
b[4240] == 4240 && 
b[4241] == 4241 && 
b[4242] == 4242 && 
b[4243] == 4243 && 
b[4244] == 4244 && 
b[4245] == 4245 && 
b[4246] == 4246 && 
b[4247] == 4247 && 
b[4248] == 4248 && 
b[4249] == 4249 && 
b[4250] == 4250 && 
b[4251] == 4251 && 
b[4252] == 4252 && 
b[4253] == 4253 && 
b[4254] == 4254 && 
b[4255] == 4255 && 
b[4256] == 4256 && 
b[4257] == 4257 && 
b[4258] == 4258 && 
b[4259] == 4259 && 
b[4260] == 4260 && 
b[4261] == 4261 && 
b[4262] == 4262 && 
b[4263] == 4263 && 
b[4264] == 4264 && 
b[4265] == 4265 && 
b[4266] == 4266 && 
b[4267] == 4267 && 
b[4268] == 4268 && 
b[4269] == 4269 && 
b[4270] == 4270 && 
b[4271] == 4271 && 
b[4272] == 4272 && 
b[4273] == 4273 && 
b[4274] == 4274 && 
b[4275] == 4275 && 
b[4276] == 4276 && 
b[4277] == 4277 && 
b[4278] == 4278 && 
b[4279] == 4279 && 
b[4280] == 4280 && 
b[4281] == 4281 && 
b[4282] == 4282 && 
b[4283] == 4283 && 
b[4284] == 4284 && 
b[4285] == 4285 && 
b[4286] == 4286 && 
b[4287] == 4287 && 
b[4288] == 4288 && 
b[4289] == 4289 && 
b[4290] == 4290 && 
b[4291] == 4291 && 
b[4292] == 4292 && 
b[4293] == 4293 && 
b[4294] == 4294 && 
b[4295] == 4295 && 
b[4296] == 4296 && 
b[4297] == 4297 && 
b[4298] == 4298 && 
b[4299] == 4299 && 
b[4300] == 4300 && 
b[4301] == 4301 && 
b[4302] == 4302 && 
b[4303] == 4303 && 
b[4304] == 4304 && 
b[4305] == 4305 && 
b[4306] == 4306 && 
b[4307] == 4307 && 
b[4308] == 4308 && 
b[4309] == 4309 && 
b[4310] == 4310 && 
b[4311] == 4311 && 
b[4312] == 4312 && 
b[4313] == 4313 && 
b[4314] == 4314 && 
b[4315] == 4315 && 
b[4316] == 4316 && 
b[4317] == 4317 && 
b[4318] == 4318 && 
b[4319] == 4319 && 
b[4320] == 4320 && 
b[4321] == 4321 && 
b[4322] == 4322 && 
b[4323] == 4323 && 
b[4324] == 4324 && 
b[4325] == 4325 && 
b[4326] == 4326 && 
b[4327] == 4327 && 
b[4328] == 4328 && 
b[4329] == 4329 && 
b[4330] == 4330 && 
b[4331] == 4331 && 
b[4332] == 4332 && 
b[4333] == 4333 && 
b[4334] == 4334 && 
b[4335] == 4335 && 
b[4336] == 4336 && 
b[4337] == 4337 && 
b[4338] == 4338 && 
b[4339] == 4339 && 
b[4340] == 4340 && 
b[4341] == 4341 && 
b[4342] == 4342 && 
b[4343] == 4343 && 
b[4344] == 4344 && 
b[4345] == 4345 && 
b[4346] == 4346 && 
b[4347] == 4347 && 
b[4348] == 4348 && 
b[4349] == 4349 && 
b[4350] == 4350 && 
b[4351] == 4351 && 
b[4352] == 4352 && 
b[4353] == 4353 && 
b[4354] == 4354 && 
b[4355] == 4355 && 
b[4356] == 4356 && 
b[4357] == 4357 && 
b[4358] == 4358 && 
b[4359] == 4359 && 
b[4360] == 4360 && 
b[4361] == 4361 && 
b[4362] == 4362 && 
b[4363] == 4363 && 
b[4364] == 4364 && 
b[4365] == 4365 && 
b[4366] == 4366 && 
b[4367] == 4367 && 
b[4368] == 4368 && 
b[4369] == 4369 && 
b[4370] == 4370 && 
b[4371] == 4371 && 
b[4372] == 4372 && 
b[4373] == 4373 && 
b[4374] == 4374 && 
b[4375] == 4375 && 
b[4376] == 4376 && 
b[4377] == 4377 && 
b[4378] == 4378 && 
b[4379] == 4379 && 
b[4380] == 4380 && 
b[4381] == 4381 && 
b[4382] == 4382 && 
b[4383] == 4383 && 
b[4384] == 4384 && 
b[4385] == 4385 && 
b[4386] == 4386 && 
b[4387] == 4387 && 
b[4388] == 4388 && 
b[4389] == 4389 && 
b[4390] == 4390 && 
b[4391] == 4391 && 
b[4392] == 4392 && 
b[4393] == 4393 && 
b[4394] == 4394 && 
b[4395] == 4395 && 
b[4396] == 4396 && 
b[4397] == 4397 && 
b[4398] == 4398 && 
b[4399] == 4399 && 
b[4400] == 4400 && 
b[4401] == 4401 && 
b[4402] == 4402 && 
b[4403] == 4403 && 
b[4404] == 4404 && 
b[4405] == 4405 && 
b[4406] == 4406 && 
b[4407] == 4407 && 
b[4408] == 4408 && 
b[4409] == 4409 && 
b[4410] == 4410 && 
b[4411] == 4411 && 
b[4412] == 4412 && 
b[4413] == 4413 && 
b[4414] == 4414 && 
b[4415] == 4415 && 
b[4416] == 4416 && 
b[4417] == 4417 && 
b[4418] == 4418 && 
b[4419] == 4419 && 
b[4420] == 4420 && 
b[4421] == 4421 && 
b[4422] == 4422 && 
b[4423] == 4423 && 
b[4424] == 4424 && 
b[4425] == 4425 && 
b[4426] == 4426 && 
b[4427] == 4427 && 
b[4428] == 4428 && 
b[4429] == 4429 && 
b[4430] == 4430 && 
b[4431] == 4431 && 
b[4432] == 4432 && 
b[4433] == 4433 && 
b[4434] == 4434 && 
b[4435] == 4435 && 
b[4436] == 4436 && 
b[4437] == 4437 && 
b[4438] == 4438 && 
b[4439] == 4439 && 
b[4440] == 4440 && 
b[4441] == 4441 && 
b[4442] == 4442 && 
b[4443] == 4443 && 
b[4444] == 4444 && 
b[4445] == 4445 && 
b[4446] == 4446 && 
b[4447] == 4447 && 
b[4448] == 4448 && 
b[4449] == 4449 && 
b[4450] == 4450 && 
b[4451] == 4451 && 
b[4452] == 4452 && 
b[4453] == 4453 && 
b[4454] == 4454 && 
b[4455] == 4455 && 
b[4456] == 4456 && 
b[4457] == 4457 && 
b[4458] == 4458 && 
b[4459] == 4459 && 
b[4460] == 4460 && 
b[4461] == 4461 && 
b[4462] == 4462 && 
b[4463] == 4463 && 
b[4464] == 4464 && 
b[4465] == 4465 && 
b[4466] == 4466 && 
b[4467] == 4467 && 
b[4468] == 4468 && 
b[4469] == 4469 && 
b[4470] == 4470 && 
b[4471] == 4471 && 
b[4472] == 4472 && 
b[4473] == 4473 && 
b[4474] == 4474 && 
b[4475] == 4475 && 
b[4476] == 4476 && 
b[4477] == 4477 && 
b[4478] == 4478 && 
b[4479] == 4479 && 
b[4480] == 4480 && 
b[4481] == 4481 && 
b[4482] == 4482 && 
b[4483] == 4483 && 
b[4484] == 4484 && 
b[4485] == 4485 && 
b[4486] == 4486 && 
b[4487] == 4487 && 
b[4488] == 4488 && 
b[4489] == 4489 && 
b[4490] == 4490 && 
b[4491] == 4491 && 
b[4492] == 4492 && 
b[4493] == 4493 && 
b[4494] == 4494 && 
b[4495] == 4495 && 
b[4496] == 4496 && 
b[4497] == 4497 && 
b[4498] == 4498 && 
b[4499] == 4499 && 
b[4500] == 4500 && 
b[4501] == 4501 && 
b[4502] == 4502 && 
b[4503] == 4503 && 
b[4504] == 4504 && 
b[4505] == 4505 && 
b[4506] == 4506 && 
b[4507] == 4507 && 
b[4508] == 4508 && 
b[4509] == 4509 && 
b[4510] == 4510 && 
b[4511] == 4511 && 
b[4512] == 4512 && 
b[4513] == 4513 && 
b[4514] == 4514 && 
b[4515] == 4515 && 
b[4516] == 4516 && 
b[4517] == 4517 && 
b[4518] == 4518 && 
b[4519] == 4519 && 
b[4520] == 4520 && 
b[4521] == 4521 && 
b[4522] == 4522 && 
b[4523] == 4523 && 
b[4524] == 4524 && 
b[4525] == 4525 && 
b[4526] == 4526 && 
b[4527] == 4527 && 
b[4528] == 4528 && 
b[4529] == 4529 && 
b[4530] == 4530 && 
b[4531] == 4531 && 
b[4532] == 4532 && 
b[4533] == 4533 && 
b[4534] == 4534 && 
b[4535] == 4535 && 
b[4536] == 4536 && 
b[4537] == 4537 && 
b[4538] == 4538 && 
b[4539] == 4539 && 
b[4540] == 4540 && 
b[4541] == 4541 && 
b[4542] == 4542 && 
b[4543] == 4543 && 
b[4544] == 4544 && 
b[4545] == 4545 && 
b[4546] == 4546 && 
b[4547] == 4547 && 
b[4548] == 4548 && 
b[4549] == 4549 && 
b[4550] == 4550 && 
b[4551] == 4551 && 
b[4552] == 4552 && 
b[4553] == 4553 && 
b[4554] == 4554 && 
b[4555] == 4555 && 
b[4556] == 4556 && 
b[4557] == 4557 && 
b[4558] == 4558 && 
b[4559] == 4559 && 
b[4560] == 4560 && 
b[4561] == 4561 && 
b[4562] == 4562 && 
b[4563] == 4563 && 
b[4564] == 4564 && 
b[4565] == 4565 && 
b[4566] == 4566 && 
b[4567] == 4567 && 
b[4568] == 4568 && 
b[4569] == 4569 && 
b[4570] == 4570 && 
b[4571] == 4571 && 
b[4572] == 4572 && 
b[4573] == 4573 && 
b[4574] == 4574 && 
b[4575] == 4575 && 
b[4576] == 4576 && 
b[4577] == 4577 && 
b[4578] == 4578 && 
b[4579] == 4579 && 
b[4580] == 4580 && 
b[4581] == 4581 && 
b[4582] == 4582 && 
b[4583] == 4583 && 
b[4584] == 4584 && 
b[4585] == 4585 && 
b[4586] == 4586 && 
b[4587] == 4587 && 
b[4588] == 4588 && 
b[4589] == 4589 && 
b[4590] == 4590 && 
b[4591] == 4591 && 
b[4592] == 4592 && 
b[4593] == 4593 && 
b[4594] == 4594 && 
b[4595] == 4595 && 
b[4596] == 4596 && 
b[4597] == 4597 && 
b[4598] == 4598 && 
b[4599] == 4599 && 
b[4600] == 4600 && 
b[4601] == 4601 && 
b[4602] == 4602 && 
b[4603] == 4603 && 
b[4604] == 4604 && 
b[4605] == 4605 && 
b[4606] == 4606 && 
b[4607] == 4607 && 
b[4608] == 4608 && 
b[4609] == 4609 && 
b[4610] == 4610 && 
b[4611] == 4611 && 
b[4612] == 4612 && 
b[4613] == 4613 && 
b[4614] == 4614 && 
b[4615] == 4615 && 
b[4616] == 4616 && 
b[4617] == 4617 && 
b[4618] == 4618 && 
b[4619] == 4619 && 
b[4620] == 4620 && 
b[4621] == 4621 && 
b[4622] == 4622 && 
b[4623] == 4623 && 
b[4624] == 4624 && 
b[4625] == 4625 && 
b[4626] == 4626 && 
b[4627] == 4627 && 
b[4628] == 4628 && 
b[4629] == 4629 && 
b[4630] == 4630 && 
b[4631] == 4631 && 
b[4632] == 4632 && 
b[4633] == 4633 && 
b[4634] == 4634 && 
b[4635] == 4635 && 
b[4636] == 4636 && 
b[4637] == 4637 && 
b[4638] == 4638 && 
b[4639] == 4639 && 
b[4640] == 4640 && 
b[4641] == 4641 && 
b[4642] == 4642 && 
b[4643] == 4643 && 
b[4644] == 4644 && 
b[4645] == 4645 && 
b[4646] == 4646 && 
b[4647] == 4647 && 
b[4648] == 4648 && 
b[4649] == 4649 && 
b[4650] == 4650 && 
b[4651] == 4651 && 
b[4652] == 4652 && 
b[4653] == 4653 && 
b[4654] == 4654 && 
b[4655] == 4655 && 
b[4656] == 4656 && 
b[4657] == 4657 && 
b[4658] == 4658 && 
b[4659] == 4659 && 
b[4660] == 4660 && 
b[4661] == 4661 && 
b[4662] == 4662 && 
b[4663] == 4663 && 
b[4664] == 4664 && 
b[4665] == 4665 && 
b[4666] == 4666 && 
b[4667] == 4667 && 
b[4668] == 4668 && 
b[4669] == 4669 && 
b[4670] == 4670 && 
b[4671] == 4671 && 
b[4672] == 4672 && 
b[4673] == 4673 && 
b[4674] == 4674 && 
b[4675] == 4675 && 
b[4676] == 4676 && 
b[4677] == 4677 && 
b[4678] == 4678 && 
b[4679] == 4679 && 
b[4680] == 4680 && 
b[4681] == 4681 && 
b[4682] == 4682 && 
b[4683] == 4683 && 
b[4684] == 4684 && 
b[4685] == 4685 && 
b[4686] == 4686 && 
b[4687] == 4687 && 
b[4688] == 4688 && 
b[4689] == 4689 && 
b[4690] == 4690 && 
b[4691] == 4691 && 
b[4692] == 4692 && 
b[4693] == 4693 && 
b[4694] == 4694 && 
b[4695] == 4695 && 
b[4696] == 4696 && 
b[4697] == 4697 && 
b[4698] == 4698 && 
b[4699] == 4699 && 
b[4700] == 4700 && 
b[4701] == 4701 && 
b[4702] == 4702 && 
b[4703] == 4703 && 
b[4704] == 4704 && 
b[4705] == 4705 && 
b[4706] == 4706 && 
b[4707] == 4707 && 
b[4708] == 4708 && 
b[4709] == 4709 && 
b[4710] == 4710 && 
b[4711] == 4711 && 
b[4712] == 4712 && 
b[4713] == 4713 && 
b[4714] == 4714 && 
b[4715] == 4715 && 
b[4716] == 4716 && 
b[4717] == 4717 && 
b[4718] == 4718 && 
b[4719] == 4719 && 
b[4720] == 4720 && 
b[4721] == 4721 && 
b[4722] == 4722 && 
b[4723] == 4723 && 
b[4724] == 4724 && 
b[4725] == 4725 && 
b[4726] == 4726 && 
b[4727] == 4727 && 
b[4728] == 4728 && 
b[4729] == 4729 && 
b[4730] == 4730 && 
b[4731] == 4731 && 
b[4732] == 4732 && 
b[4733] == 4733 && 
b[4734] == 4734 && 
b[4735] == 4735 && 
b[4736] == 4736 && 
b[4737] == 4737 && 
b[4738] == 4738 && 
b[4739] == 4739 && 
b[4740] == 4740 && 
b[4741] == 4741 && 
b[4742] == 4742 && 
b[4743] == 4743 && 
b[4744] == 4744 && 
b[4745] == 4745 && 
b[4746] == 4746 && 
b[4747] == 4747 && 
b[4748] == 4748 && 
b[4749] == 4749 && 
b[4750] == 4750 && 
b[4751] == 4751 && 
b[4752] == 4752 && 
b[4753] == 4753 && 
b[4754] == 4754 && 
b[4755] == 4755 && 
b[4756] == 4756 && 
b[4757] == 4757 && 
b[4758] == 4758 && 
b[4759] == 4759 && 
b[4760] == 4760 && 
b[4761] == 4761 && 
b[4762] == 4762 && 
b[4763] == 4763 && 
b[4764] == 4764 && 
b[4765] == 4765 && 
b[4766] == 4766 && 
b[4767] == 4767 && 
b[4768] == 4768 && 
b[4769] == 4769 && 
b[4770] == 4770 && 
b[4771] == 4771 && 
b[4772] == 4772 && 
b[4773] == 4773 && 
b[4774] == 4774 && 
b[4775] == 4775 && 
b[4776] == 4776 && 
b[4777] == 4777 && 
b[4778] == 4778 && 
b[4779] == 4779 && 
b[4780] == 4780 && 
b[4781] == 4781 && 
b[4782] == 4782 && 
b[4783] == 4783 && 
b[4784] == 4784 && 
b[4785] == 4785 && 
b[4786] == 4786 && 
b[4787] == 4787 && 
b[4788] == 4788 && 
b[4789] == 4789 && 
b[4790] == 4790 && 
b[4791] == 4791 && 
b[4792] == 4792 && 
b[4793] == 4793 && 
b[4794] == 4794 && 
b[4795] == 4795 && 
b[4796] == 4796 && 
b[4797] == 4797 && 
b[4798] == 4798 && 
b[4799] == 4799 && 
b[4800] == 4800 && 
b[4801] == 4801 && 
b[4802] == 4802 && 
b[4803] == 4803 && 
b[4804] == 4804 && 
b[4805] == 4805 && 
b[4806] == 4806 && 
b[4807] == 4807 && 
b[4808] == 4808 && 
b[4809] == 4809 && 
b[4810] == 4810 && 
b[4811] == 4811 && 
b[4812] == 4812 && 
b[4813] == 4813 && 
b[4814] == 4814 && 
b[4815] == 4815 && 
b[4816] == 4816 && 
b[4817] == 4817 && 
b[4818] == 4818 && 
b[4819] == 4819 && 
b[4820] == 4820 && 
b[4821] == 4821 && 
b[4822] == 4822 && 
b[4823] == 4823 && 
b[4824] == 4824 && 
b[4825] == 4825 && 
b[4826] == 4826 && 
b[4827] == 4827 && 
b[4828] == 4828 && 
b[4829] == 4829 && 
b[4830] == 4830 && 
b[4831] == 4831 && 
b[4832] == 4832 && 
b[4833] == 4833 && 
b[4834] == 4834 && 
b[4835] == 4835 && 
b[4836] == 4836 && 
b[4837] == 4837 && 
b[4838] == 4838 && 
b[4839] == 4839 && 
b[4840] == 4840 && 
b[4841] == 4841 && 
b[4842] == 4842 && 
b[4843] == 4843 && 
b[4844] == 4844 && 
b[4845] == 4845 && 
b[4846] == 4846 && 
b[4847] == 4847 && 
b[4848] == 4848 && 
b[4849] == 4849 && 
b[4850] == 4850 && 
b[4851] == 4851 && 
b[4852] == 4852 && 
b[4853] == 4853 && 
b[4854] == 4854 && 
b[4855] == 4855 && 
b[4856] == 4856 && 
b[4857] == 4857 && 
b[4858] == 4858 && 
b[4859] == 4859 && 
b[4860] == 4860 && 
b[4861] == 4861 && 
b[4862] == 4862 && 
b[4863] == 4863 && 
b[4864] == 4864 && 
b[4865] == 4865 && 
b[4866] == 4866 && 
b[4867] == 4867 && 
b[4868] == 4868 && 
b[4869] == 4869 && 
b[4870] == 4870 && 
b[4871] == 4871 && 
b[4872] == 4872 && 
b[4873] == 4873 && 
b[4874] == 4874 && 
b[4875] == 4875 && 
b[4876] == 4876 && 
b[4877] == 4877 && 
b[4878] == 4878 && 
b[4879] == 4879 && 
b[4880] == 4880 && 
b[4881] == 4881 && 
b[4882] == 4882 && 
b[4883] == 4883 && 
b[4884] == 4884 && 
b[4885] == 4885 && 
b[4886] == 4886 && 
b[4887] == 4887 && 
b[4888] == 4888 && 
b[4889] == 4889 && 
b[4890] == 4890 && 
b[4891] == 4891 && 
b[4892] == 4892 && 
b[4893] == 4893 && 
b[4894] == 4894 && 
b[4895] == 4895 && 
b[4896] == 4896 && 
b[4897] == 4897 && 
b[4898] == 4898 && 
b[4899] == 4899 && 
b[4900] == 4900 && 
b[4901] == 4901 && 
b[4902] == 4902 && 
b[4903] == 4903 && 
b[4904] == 4904 && 
b[4905] == 4905 && 
b[4906] == 4906 && 
b[4907] == 4907 && 
b[4908] == 4908 && 
b[4909] == 4909 && 
b[4910] == 4910 && 
b[4911] == 4911 && 
b[4912] == 4912 && 
b[4913] == 4913 && 
b[4914] == 4914 && 
b[4915] == 4915 && 
b[4916] == 4916 && 
b[4917] == 4917 && 
b[4918] == 4918 && 
b[4919] == 4919 && 
b[4920] == 4920 && 
b[4921] == 4921 && 
b[4922] == 4922 && 
b[4923] == 4923 && 
b[4924] == 4924 && 
b[4925] == 4925 && 
b[4926] == 4926 && 
b[4927] == 4927 && 
b[4928] == 4928 && 
b[4929] == 4929 && 
b[4930] == 4930 && 
b[4931] == 4931 && 
b[4932] == 4932 && 
b[4933] == 4933 && 
b[4934] == 4934 && 
b[4935] == 4935 && 
b[4936] == 4936 && 
b[4937] == 4937 && 
b[4938] == 4938 && 
b[4939] == 4939 && 
b[4940] == 4940 && 
b[4941] == 4941 && 
b[4942] == 4942 && 
b[4943] == 4943 && 
b[4944] == 4944 && 
b[4945] == 4945 && 
b[4946] == 4946 && 
b[4947] == 4947 && 
b[4948] == 4948 && 
b[4949] == 4949 && 
b[4950] == 4950 && 
b[4951] == 4951 && 
b[4952] == 4952 && 
b[4953] == 4953 && 
b[4954] == 4954 && 
b[4955] == 4955 && 
b[4956] == 4956 && 
b[4957] == 4957 && 
b[4958] == 4958 && 
b[4959] == 4959 && 
b[4960] == 4960 && 
b[4961] == 4961 && 
b[4962] == 4962 && 
b[4963] == 4963 && 
b[4964] == 4964 && 
b[4965] == 4965 && 
b[4966] == 4966 && 
b[4967] == 4967 && 
b[4968] == 4968 && 
b[4969] == 4969 && 
b[4970] == 4970 && 
b[4971] == 4971 && 
b[4972] == 4972 && 
b[4973] == 4973 && 
b[4974] == 4974 && 
b[4975] == 4975 && 
b[4976] == 4976 && 
b[4977] == 4977 && 
b[4978] == 4978 && 
b[4979] == 4979 && 
b[4980] == 4980 && 
b[4981] == 4981 && 
b[4982] == 4982 && 
b[4983] == 4983 && 
b[4984] == 4984 && 
b[4985] == 4985 && 
b[4986] == 4986 && 
b[4987] == 4987 && 
b[4988] == 4988 && 
b[4989] == 4989 && 
b[4990] == 4990 && 
b[4991] == 4991 && 
b[4992] == 4992 && 
b[4993] == 4993 && 
b[4994] == 4994 && 
b[4995] == 4995 && 
b[4996] == 4996 && 
b[4997] == 4997 && 
b[4998] == 4998 && 
b[4999] == 4999 && 
b[5000] == 5000 && 
b[5001] == 5001 && 
b[5002] == 5002 && 
b[5003] == 5003 && 
b[5004] == 5004 && 
b[5005] == 5005 && 
b[5006] == 5006 && 
b[5007] == 5007 && 
b[5008] == 5008 && 
b[5009] == 5009 && 
b[5010] == 5010 && 
b[5011] == 5011 && 
b[5012] == 5012 && 
b[5013] == 5013 && 
b[5014] == 5014 && 
b[5015] == 5015 && 
b[5016] == 5016 && 
b[5017] == 5017 && 
b[5018] == 5018 && 
b[5019] == 5019 && 
b[5020] == 5020 && 
b[5021] == 5021 && 
b[5022] == 5022 && 
b[5023] == 5023 && 
b[5024] == 5024 && 
b[5025] == 5025 && 
b[5026] == 5026 && 
b[5027] == 5027 && 
b[5028] == 5028 && 
b[5029] == 5029 && 
b[5030] == 5030 && 
b[5031] == 5031 && 
b[5032] == 5032 && 
b[5033] == 5033 && 
b[5034] == 5034 && 
b[5035] == 5035 && 
b[5036] == 5036 && 
b[5037] == 5037 && 
b[5038] == 5038 && 
b[5039] == 5039 && 
b[5040] == 5040 && 
b[5041] == 5041 && 
b[5042] == 5042 && 
b[5043] == 5043 && 
b[5044] == 5044 && 
b[5045] == 5045 && 
b[5046] == 5046 && 
b[5047] == 5047 && 
b[5048] == 5048 && 
b[5049] == 5049 && 
b[5050] == 5050 && 
b[5051] == 5051 && 
b[5052] == 5052 && 
b[5053] == 5053 && 
b[5054] == 5054 && 
b[5055] == 5055 && 
b[5056] == 5056 && 
b[5057] == 5057 && 
b[5058] == 5058 && 
b[5059] == 5059 && 
b[5060] == 5060 && 
b[5061] == 5061 && 
b[5062] == 5062 && 
b[5063] == 5063 && 
b[5064] == 5064 && 
b[5065] == 5065 && 
b[5066] == 5066 && 
b[5067] == 5067 && 
b[5068] == 5068 && 
b[5069] == 5069 && 
b[5070] == 5070 && 
b[5071] == 5071 && 
b[5072] == 5072 && 
b[5073] == 5073 && 
b[5074] == 5074 && 
b[5075] == 5075 && 
b[5076] == 5076 && 
b[5077] == 5077 && 
b[5078] == 5078 && 
b[5079] == 5079 && 
b[5080] == 5080 && 
b[5081] == 5081 && 
b[5082] == 5082 && 
b[5083] == 5083 && 
b[5084] == 5084 && 
b[5085] == 5085 && 
b[5086] == 5086 && 
b[5087] == 5087 && 
b[5088] == 5088 && 
b[5089] == 5089 && 
b[5090] == 5090 && 
b[5091] == 5091 && 
b[5092] == 5092 && 
b[5093] == 5093 && 
b[5094] == 5094 && 
b[5095] == 5095 && 
b[5096] == 5096 && 
b[5097] == 5097 && 
b[5098] == 5098 && 
b[5099] == 5099 && 
b[5100] == 5100 && 
b[5101] == 5101 && 
b[5102] == 5102 && 
b[5103] == 5103 && 
b[5104] == 5104 && 
b[5105] == 5105 && 
b[5106] == 5106 && 
b[5107] == 5107 && 
b[5108] == 5108 && 
b[5109] == 5109 && 
b[5110] == 5110 && 
b[5111] == 5111 && 
b[5112] == 5112 && 
b[5113] == 5113 && 
b[5114] == 5114 && 
b[5115] == 5115 && 
b[5116] == 5116 && 
b[5117] == 5117 && 
b[5118] == 5118 && 
b[5119] == 5119 && 
b[5120] == 5120 && 
b[5121] == 5121 && 
b[5122] == 5122 && 
b[5123] == 5123 && 
b[5124] == 5124 && 
b[5125] == 5125 && 
b[5126] == 5126 && 
b[5127] == 5127 && 
b[5128] == 5128 && 
b[5129] == 5129 && 
b[5130] == 5130 && 
b[5131] == 5131 && 
b[5132] == 5132 && 
b[5133] == 5133 && 
b[5134] == 5134 && 
b[5135] == 5135 && 
b[5136] == 5136 && 
b[5137] == 5137 && 
b[5138] == 5138 && 
b[5139] == 5139 && 
b[5140] == 5140 && 
b[5141] == 5141 && 
b[5142] == 5142 && 
b[5143] == 5143 && 
b[5144] == 5144 && 
b[5145] == 5145 && 
b[5146] == 5146 && 
b[5147] == 5147 && 
b[5148] == 5148 && 
b[5149] == 5149 && 
b[5150] == 5150 && 
b[5151] == 5151 && 
b[5152] == 5152 && 
b[5153] == 5153 && 
b[5154] == 5154 && 
b[5155] == 5155 && 
b[5156] == 5156 && 
b[5157] == 5157 && 
b[5158] == 5158 && 
b[5159] == 5159 && 
b[5160] == 5160 && 
b[5161] == 5161 && 
b[5162] == 5162 && 
b[5163] == 5163 && 
b[5164] == 5164 && 
b[5165] == 5165 && 
b[5166] == 5166 && 
b[5167] == 5167 && 
b[5168] == 5168 && 
b[5169] == 5169 && 
b[5170] == 5170 && 
b[5171] == 5171 && 
b[5172] == 5172 && 
b[5173] == 5173 && 
b[5174] == 5174 && 
b[5175] == 5175 && 
b[5176] == 5176 && 
b[5177] == 5177 && 
b[5178] == 5178 && 
b[5179] == 5179 && 
b[5180] == 5180 && 
b[5181] == 5181 && 
b[5182] == 5182 && 
b[5183] == 5183 && 
b[5184] == 5184 && 
b[5185] == 5185 && 
b[5186] == 5186 && 
b[5187] == 5187 && 
b[5188] == 5188 && 
b[5189] == 5189 && 
b[5190] == 5190 && 
b[5191] == 5191 && 
b[5192] == 5192 && 
b[5193] == 5193 && 
b[5194] == 5194 && 
b[5195] == 5195 && 
b[5196] == 5196 && 
b[5197] == 5197 && 
b[5198] == 5198 && 
b[5199] == 5199 && 
b[5200] == 5200 && 
b[5201] == 5201 && 
b[5202] == 5202 && 
b[5203] == 5203 && 
b[5204] == 5204 && 
b[5205] == 5205 && 
b[5206] == 5206 && 
b[5207] == 5207 && 
b[5208] == 5208 && 
b[5209] == 5209 && 
b[5210] == 5210 && 
b[5211] == 5211 && 
b[5212] == 5212 && 
b[5213] == 5213 && 
b[5214] == 5214 && 
b[5215] == 5215 && 
b[5216] == 5216 && 
b[5217] == 5217 && 
b[5218] == 5218 && 
b[5219] == 5219 && 
b[5220] == 5220 && 
b[5221] == 5221 && 
b[5222] == 5222 && 
b[5223] == 5223 && 
b[5224] == 5224 && 
b[5225] == 5225 && 
b[5226] == 5226 && 
b[5227] == 5227 && 
b[5228] == 5228 && 
b[5229] == 5229 && 
b[5230] == 5230 && 
b[5231] == 5231 && 
b[5232] == 5232 && 
b[5233] == 5233 && 
b[5234] == 5234 && 
b[5235] == 5235 && 
b[5236] == 5236 && 
b[5237] == 5237 && 
b[5238] == 5238 && 
b[5239] == 5239 && 
b[5240] == 5240 && 
b[5241] == 5241 && 
b[5242] == 5242 && 
b[5243] == 5243 && 
b[5244] == 5244 && 
b[5245] == 5245 && 
b[5246] == 5246 && 
b[5247] == 5247 && 
b[5248] == 5248 && 
b[5249] == 5249 && 
b[5250] == 5250 && 
b[5251] == 5251 && 
b[5252] == 5252 && 
b[5253] == 5253 && 
b[5254] == 5254 && 
b[5255] == 5255 && 
b[5256] == 5256 && 
b[5257] == 5257 && 
b[5258] == 5258 && 
b[5259] == 5259 && 
b[5260] == 5260 && 
b[5261] == 5261 && 
b[5262] == 5262 && 
b[5263] == 5263 && 
b[5264] == 5264 && 
b[5265] == 5265 && 
b[5266] == 5266 && 
b[5267] == 5267 && 
b[5268] == 5268 && 
b[5269] == 5269 && 
b[5270] == 5270 && 
b[5271] == 5271 && 
b[5272] == 5272 && 
b[5273] == 5273 && 
b[5274] == 5274 && 
b[5275] == 5275 && 
b[5276] == 5276 && 
b[5277] == 5277 && 
b[5278] == 5278 && 
b[5279] == 5279 && 
b[5280] == 5280 && 
b[5281] == 5281 && 
b[5282] == 5282 && 
b[5283] == 5283 && 
b[5284] == 5284 && 
b[5285] == 5285 && 
b[5286] == 5286 && 
b[5287] == 5287 && 
b[5288] == 5288 && 
b[5289] == 5289 && 
b[5290] == 5290 && 
b[5291] == 5291 && 
b[5292] == 5292 && 
b[5293] == 5293 && 
b[5294] == 5294 && 
b[5295] == 5295 && 
b[5296] == 5296 && 
b[5297] == 5297 && 
b[5298] == 5298 && 
b[5299] == 5299 && 
b[5300] == 5300 && 
b[5301] == 5301 && 
b[5302] == 5302 && 
b[5303] == 5303 && 
b[5304] == 5304 && 
b[5305] == 5305 && 
b[5306] == 5306 && 
b[5307] == 5307 && 
b[5308] == 5308 && 
b[5309] == 5309 && 
b[5310] == 5310 && 
b[5311] == 5311 && 
b[5312] == 5312 && 
b[5313] == 5313 && 
b[5314] == 5314 && 
b[5315] == 5315 && 
b[5316] == 5316 && 
b[5317] == 5317 && 
b[5318] == 5318 && 
b[5319] == 5319 && 
b[5320] == 5320 && 
b[5321] == 5321 && 
b[5322] == 5322 && 
b[5323] == 5323 && 
b[5324] == 5324 && 
b[5325] == 5325 && 
b[5326] == 5326 && 
b[5327] == 5327 && 
b[5328] == 5328 && 
b[5329] == 5329 && 
b[5330] == 5330 && 
b[5331] == 5331 && 
b[5332] == 5332 && 
b[5333] == 5333 && 
b[5334] == 5334 && 
b[5335] == 5335 && 
b[5336] == 5336 && 
b[5337] == 5337 && 
b[5338] == 5338 && 
b[5339] == 5339 && 
b[5340] == 5340 && 
b[5341] == 5341 && 
b[5342] == 5342 && 
b[5343] == 5343 && 
b[5344] == 5344 && 
b[5345] == 5345 && 
b[5346] == 5346 && 
b[5347] == 5347 && 
b[5348] == 5348 && 
b[5349] == 5349 && 
b[5350] == 5350 && 
b[5351] == 5351 && 
b[5352] == 5352 && 
b[5353] == 5353 && 
b[5354] == 5354 && 
b[5355] == 5355 && 
b[5356] == 5356 && 
b[5357] == 5357 && 
b[5358] == 5358 && 
b[5359] == 5359 && 
b[5360] == 5360 && 
b[5361] == 5361 && 
b[5362] == 5362 && 
b[5363] == 5363 && 
b[5364] == 5364 && 
b[5365] == 5365 && 
b[5366] == 5366 && 
b[5367] == 5367 && 
b[5368] == 5368 && 
b[5369] == 5369 && 
b[5370] == 5370 && 
b[5371] == 5371 && 
b[5372] == 5372 && 
b[5373] == 5373 && 
b[5374] == 5374 && 
b[5375] == 5375 && 
b[5376] == 5376 && 
b[5377] == 5377 && 
b[5378] == 5378 && 
b[5379] == 5379 && 
b[5380] == 5380 && 
b[5381] == 5381 && 
b[5382] == 5382 && 
b[5383] == 5383 && 
b[5384] == 5384 && 
b[5385] == 5385 && 
b[5386] == 5386 && 
b[5387] == 5387 && 
b[5388] == 5388 && 
b[5389] == 5389 && 
b[5390] == 5390 && 
b[5391] == 5391 && 
b[5392] == 5392 && 
b[5393] == 5393 && 
b[5394] == 5394 && 
b[5395] == 5395 && 
b[5396] == 5396 && 
b[5397] == 5397 && 
b[5398] == 5398 && 
b[5399] == 5399 && 
b[5400] == 5400 && 
b[5401] == 5401 && 
b[5402] == 5402 && 
b[5403] == 5403 && 
b[5404] == 5404 && 
b[5405] == 5405 && 
b[5406] == 5406 && 
b[5407] == 5407 && 
b[5408] == 5408 && 
b[5409] == 5409 && 
b[5410] == 5410 && 
b[5411] == 5411 && 
b[5412] == 5412 && 
b[5413] == 5413 && 
b[5414] == 5414 && 
b[5415] == 5415 && 
b[5416] == 5416 && 
b[5417] == 5417 && 
b[5418] == 5418 && 
b[5419] == 5419 && 
b[5420] == 5420 && 
b[5421] == 5421 && 
b[5422] == 5422 && 
b[5423] == 5423 && 
b[5424] == 5424 && 
b[5425] == 5425 && 
b[5426] == 5426 && 
b[5427] == 5427 && 
b[5428] == 5428 && 
b[5429] == 5429 && 
b[5430] == 5430 && 
b[5431] == 5431 && 
b[5432] == 5432 && 
b[5433] == 5433 && 
b[5434] == 5434 && 
b[5435] == 5435 && 
b[5436] == 5436 && 
b[5437] == 5437 && 
b[5438] == 5438 && 
b[5439] == 5439 && 
b[5440] == 5440 && 
b[5441] == 5441 && 
b[5442] == 5442 && 
b[5443] == 5443 && 
b[5444] == 5444 && 
b[5445] == 5445 && 
b[5446] == 5446 && 
b[5447] == 5447 && 
b[5448] == 5448 && 
b[5449] == 5449 && 
b[5450] == 5450 && 
b[5451] == 5451 && 
b[5452] == 5452 && 
b[5453] == 5453 && 
b[5454] == 5454 && 
b[5455] == 5455 && 
b[5456] == 5456 && 
b[5457] == 5457 && 
b[5458] == 5458 && 
b[5459] == 5459 && 
b[5460] == 5460 && 
b[5461] == 5461 && 
b[5462] == 5462 && 
b[5463] == 5463 && 
b[5464] == 5464 && 
b[5465] == 5465 && 
b[5466] == 5466 && 
b[5467] == 5467 && 
b[5468] == 5468 && 
b[5469] == 5469 && 
b[5470] == 5470 && 
b[5471] == 5471 && 
b[5472] == 5472 && 
b[5473] == 5473 && 
b[5474] == 5474 && 
b[5475] == 5475 && 
b[5476] == 5476 && 
b[5477] == 5477 && 
b[5478] == 5478 && 
b[5479] == 5479 && 
b[5480] == 5480 && 
b[5481] == 5481 && 
b[5482] == 5482 && 
b[5483] == 5483 && 
b[5484] == 5484 && 
b[5485] == 5485 && 
b[5486] == 5486 && 
b[5487] == 5487 && 
b[5488] == 5488 && 
b[5489] == 5489 && 
b[5490] == 5490 && 
b[5491] == 5491 && 
b[5492] == 5492 && 
b[5493] == 5493 && 
b[5494] == 5494 && 
b[5495] == 5495 && 
b[5496] == 5496 && 
b[5497] == 5497 && 
b[5498] == 5498 && 
b[5499] == 5499 && 
b[5500] == 5500 && 
b[5501] == 5501 && 
b[5502] == 5502 && 
b[5503] == 5503 && 
b[5504] == 5504 && 
b[5505] == 5505 && 
b[5506] == 5506 && 
b[5507] == 5507 && 
b[5508] == 5508 && 
b[5509] == 5509 && 
b[5510] == 5510 && 
b[5511] == 5511 && 
b[5512] == 5512 && 
b[5513] == 5513 && 
b[5514] == 5514 && 
b[5515] == 5515 && 
b[5516] == 5516 && 
b[5517] == 5517 && 
b[5518] == 5518 && 
b[5519] == 5519 && 
b[5520] == 5520 && 
b[5521] == 5521 && 
b[5522] == 5522 && 
b[5523] == 5523 && 
b[5524] == 5524 && 
b[5525] == 5525 && 
b[5526] == 5526 && 
b[5527] == 5527 && 
b[5528] == 5528 && 
b[5529] == 5529 && 
b[5530] == 5530 && 
b[5531] == 5531 && 
b[5532] == 5532 && 
b[5533] == 5533 && 
b[5534] == 5534 && 
b[5535] == 5535 && 
b[5536] == 5536 && 
b[5537] == 5537 && 
b[5538] == 5538 && 
b[5539] == 5539 && 
b[5540] == 5540 && 
b[5541] == 5541 && 
b[5542] == 5542 && 
b[5543] == 5543 && 
b[5544] == 5544 && 
b[5545] == 5545 && 
b[5546] == 5546 && 
b[5547] == 5547 && 
b[5548] == 5548 && 
b[5549] == 5549 && 
b[5550] == 5550 && 
b[5551] == 5551 && 
b[5552] == 5552 && 
b[5553] == 5553 && 
b[5554] == 5554 && 
b[5555] == 5555 && 
b[5556] == 5556 && 
b[5557] == 5557 && 
b[5558] == 5558 && 
b[5559] == 5559 && 
b[5560] == 5560 && 
b[5561] == 5561 && 
b[5562] == 5562 && 
b[5563] == 5563 && 
b[5564] == 5564 && 
b[5565] == 5565 && 
b[5566] == 5566 && 
b[5567] == 5567 && 
b[5568] == 5568 && 
b[5569] == 5569 && 
b[5570] == 5570 && 
b[5571] == 5571 && 
b[5572] == 5572 && 
b[5573] == 5573 && 
b[5574] == 5574 && 
b[5575] == 5575 && 
b[5576] == 5576 && 
b[5577] == 5577 && 
b[5578] == 5578 && 
b[5579] == 5579 && 
b[5580] == 5580 && 
b[5581] == 5581 && 
b[5582] == 5582 && 
b[5583] == 5583 && 
b[5584] == 5584 && 
b[5585] == 5585 && 
b[5586] == 5586 && 
b[5587] == 5587 && 
b[5588] == 5588 && 
b[5589] == 5589 && 
b[5590] == 5590 && 
b[5591] == 5591 && 
b[5592] == 5592 && 
b[5593] == 5593 && 
b[5594] == 5594 && 
b[5595] == 5595 && 
b[5596] == 5596 && 
b[5597] == 5597 && 
b[5598] == 5598 && 
b[5599] == 5599 && 
b[5600] == 5600 && 
b[5601] == 5601 && 
b[5602] == 5602 && 
b[5603] == 5603 && 
b[5604] == 5604 && 
b[5605] == 5605 && 
b[5606] == 5606 && 
b[5607] == 5607 && 
b[5608] == 5608 && 
b[5609] == 5609 && 
b[5610] == 5610 && 
b[5611] == 5611 && 
b[5612] == 5612 && 
b[5613] == 5613 && 
b[5614] == 5614 && 
b[5615] == 5615 && 
b[5616] == 5616 && 
b[5617] == 5617 && 
b[5618] == 5618 && 
b[5619] == 5619 && 
b[5620] == 5620 && 
b[5621] == 5621 && 
b[5622] == 5622 && 
b[5623] == 5623 && 
b[5624] == 5624 && 
b[5625] == 5625 && 
b[5626] == 5626 && 
b[5627] == 5627 && 
b[5628] == 5628 && 
b[5629] == 5629 && 
b[5630] == 5630 && 
b[5631] == 5631 && 
b[5632] == 5632 && 
b[5633] == 5633 && 
b[5634] == 5634 && 
b[5635] == 5635 && 
b[5636] == 5636 && 
b[5637] == 5637 && 
b[5638] == 5638 && 
b[5639] == 5639 && 
b[5640] == 5640 && 
b[5641] == 5641 && 
b[5642] == 5642 && 
b[5643] == 5643 && 
b[5644] == 5644 && 
b[5645] == 5645 && 
b[5646] == 5646 && 
b[5647] == 5647 && 
b[5648] == 5648 && 
b[5649] == 5649 && 
b[5650] == 5650 && 
b[5651] == 5651 && 
b[5652] == 5652 && 
b[5653] == 5653 && 
b[5654] == 5654 && 
b[5655] == 5655 && 
b[5656] == 5656 && 
b[5657] == 5657 && 
b[5658] == 5658 && 
b[5659] == 5659 && 
b[5660] == 5660 && 
b[5661] == 5661 && 
b[5662] == 5662 && 
b[5663] == 5663 && 
b[5664] == 5664 && 
b[5665] == 5665 && 
b[5666] == 5666 && 
b[5667] == 5667 && 
b[5668] == 5668 && 
b[5669] == 5669 && 
b[5670] == 5670 && 
b[5671] == 5671 && 
b[5672] == 5672 && 
b[5673] == 5673 && 
b[5674] == 5674 && 
b[5675] == 5675 && 
b[5676] == 5676 && 
b[5677] == 5677 && 
b[5678] == 5678 && 
b[5679] == 5679 && 
b[5680] == 5680 && 
b[5681] == 5681 && 
b[5682] == 5682 && 
b[5683] == 5683 && 
b[5684] == 5684 && 
b[5685] == 5685 && 
b[5686] == 5686 && 
b[5687] == 5687 && 
b[5688] == 5688 && 
b[5689] == 5689 && 
b[5690] == 5690 && 
b[5691] == 5691 && 
b[5692] == 5692 && 
b[5693] == 5693 && 
b[5694] == 5694 && 
b[5695] == 5695 && 
b[5696] == 5696 && 
b[5697] == 5697 && 
b[5698] == 5698 && 
b[5699] == 5699 && 
b[5700] == 5700 && 
b[5701] == 5701 && 
b[5702] == 5702 && 
b[5703] == 5703 && 
b[5704] == 5704 && 
b[5705] == 5705 && 
b[5706] == 5706 && 
b[5707] == 5707 && 
b[5708] == 5708 && 
b[5709] == 5709 && 
b[5710] == 5710 && 
b[5711] == 5711 && 
b[5712] == 5712 && 
b[5713] == 5713 && 
b[5714] == 5714 && 
b[5715] == 5715 && 
b[5716] == 5716 && 
b[5717] == 5717 && 
b[5718] == 5718 && 
b[5719] == 5719 && 
b[5720] == 5720 && 
b[5721] == 5721 && 
b[5722] == 5722 && 
b[5723] == 5723 && 
b[5724] == 5724 && 
b[5725] == 5725 && 
b[5726] == 5726 && 
b[5727] == 5727 && 
b[5728] == 5728 && 
b[5729] == 5729 && 
b[5730] == 5730 && 
b[5731] == 5731 && 
b[5732] == 5732 && 
b[5733] == 5733 && 
b[5734] == 5734 && 
b[5735] == 5735 && 
b[5736] == 5736 && 
b[5737] == 5737 && 
b[5738] == 5738 && 
b[5739] == 5739 && 
b[5740] == 5740 && 
b[5741] == 5741 && 
b[5742] == 5742 && 
b[5743] == 5743 && 
b[5744] == 5744 && 
b[5745] == 5745 && 
b[5746] == 5746 && 
b[5747] == 5747 && 
b[5748] == 5748 && 
b[5749] == 5749 && 
b[5750] == 5750 && 
b[5751] == 5751 && 
b[5752] == 5752 && 
b[5753] == 5753 && 
b[5754] == 5754 && 
b[5755] == 5755 && 
b[5756] == 5756 && 
b[5757] == 5757 && 
b[5758] == 5758 && 
b[5759] == 5759 && 
b[5760] == 5760 && 
b[5761] == 5761 && 
b[5762] == 5762 && 
b[5763] == 5763 && 
b[5764] == 5764 && 
b[5765] == 5765 && 
b[5766] == 5766 && 
b[5767] == 5767 && 
b[5768] == 5768 && 
b[5769] == 5769 && 
b[5770] == 5770 && 
b[5771] == 5771 && 
b[5772] == 5772 && 
b[5773] == 5773 && 
b[5774] == 5774 && 
b[5775] == 5775 && 
b[5776] == 5776 && 
b[5777] == 5777 && 
b[5778] == 5778 && 
b[5779] == 5779 && 
b[5780] == 5780 && 
b[5781] == 5781 && 
b[5782] == 5782 && 
b[5783] == 5783 && 
b[5784] == 5784 && 
b[5785] == 5785 && 
b[5786] == 5786 && 
b[5787] == 5787 && 
b[5788] == 5788 && 
b[5789] == 5789 && 
b[5790] == 5790 && 
b[5791] == 5791 && 
b[5792] == 5792 && 
b[5793] == 5793 && 
b[5794] == 5794 && 
b[5795] == 5795 && 
b[5796] == 5796 && 
b[5797] == 5797 && 
b[5798] == 5798 && 
b[5799] == 5799 && 
b[5800] == 5800 && 
b[5801] == 5801 && 
b[5802] == 5802 && 
b[5803] == 5803 && 
b[5804] == 5804 && 
b[5805] == 5805 && 
b[5806] == 5806 && 
b[5807] == 5807 && 
b[5808] == 5808 && 
b[5809] == 5809 && 
b[5810] == 5810 && 
b[5811] == 5811 && 
b[5812] == 5812 && 
b[5813] == 5813 && 
b[5814] == 5814 && 
b[5815] == 5815 && 
b[5816] == 5816 && 
b[5817] == 5817 && 
b[5818] == 5818 && 
b[5819] == 5819 && 
b[5820] == 5820 && 
b[5821] == 5821 && 
b[5822] == 5822 && 
b[5823] == 5823 && 
b[5824] == 5824 && 
b[5825] == 5825 && 
b[5826] == 5826 && 
b[5827] == 5827 && 
b[5828] == 5828 && 
b[5829] == 5829 && 
b[5830] == 5830 && 
b[5831] == 5831 && 
b[5832] == 5832 && 
b[5833] == 5833 && 
b[5834] == 5834 && 
b[5835] == 5835 && 
b[5836] == 5836 && 
b[5837] == 5837 && 
b[5838] == 5838 && 
b[5839] == 5839 && 
b[5840] == 5840 && 
b[5841] == 5841 && 
b[5842] == 5842 && 
b[5843] == 5843 && 
b[5844] == 5844 && 
b[5845] == 5845 && 
b[5846] == 5846 && 
b[5847] == 5847 && 
b[5848] == 5848 && 
b[5849] == 5849 && 
b[5850] == 5850 && 
b[5851] == 5851 && 
b[5852] == 5852 && 
b[5853] == 5853 && 
b[5854] == 5854 && 
b[5855] == 5855 && 
b[5856] == 5856 && 
b[5857] == 5857 && 
b[5858] == 5858 && 
b[5859] == 5859 && 
b[5860] == 5860 && 
b[5861] == 5861 && 
b[5862] == 5862 && 
b[5863] == 5863 && 
b[5864] == 5864 && 
b[5865] == 5865 && 
b[5866] == 5866 && 
b[5867] == 5867 && 
b[5868] == 5868 && 
b[5869] == 5869 && 
b[5870] == 5870 && 
b[5871] == 5871 && 
b[5872] == 5872 && 
b[5873] == 5873 && 
b[5874] == 5874 && 
b[5875] == 5875 && 
b[5876] == 5876 && 
b[5877] == 5877 && 
b[5878] == 5878 && 
b[5879] == 5879 && 
b[5880] == 5880 && 
b[5881] == 5881 && 
b[5882] == 5882 && 
b[5883] == 5883 && 
b[5884] == 5884 && 
b[5885] == 5885 && 
b[5886] == 5886 && 
b[5887] == 5887 && 
b[5888] == 5888 && 
b[5889] == 5889 && 
b[5890] == 5890 && 
b[5891] == 5891 && 
b[5892] == 5892 && 
b[5893] == 5893 && 
b[5894] == 5894 && 
b[5895] == 5895 && 
b[5896] == 5896 && 
b[5897] == 5897 && 
b[5898] == 5898 && 
b[5899] == 5899 && 
b[5900] == 5900 && 
b[5901] == 5901 && 
b[5902] == 5902 && 
b[5903] == 5903 && 
b[5904] == 5904 && 
b[5905] == 5905 && 
b[5906] == 5906 && 
b[5907] == 5907 && 
b[5908] == 5908 && 
b[5909] == 5909 && 
b[5910] == 5910 && 
b[5911] == 5911 && 
b[5912] == 5912 && 
b[5913] == 5913 && 
b[5914] == 5914 && 
b[5915] == 5915 && 
b[5916] == 5916 && 
b[5917] == 5917 && 
b[5918] == 5918 && 
b[5919] == 5919 && 
b[5920] == 5920 && 
b[5921] == 5921 && 
b[5922] == 5922 && 
b[5923] == 5923 && 
b[5924] == 5924 && 
b[5925] == 5925 && 
b[5926] == 5926 && 
b[5927] == 5927 && 
b[5928] == 5928 && 
b[5929] == 5929 && 
b[5930] == 5930 && 
b[5931] == 5931 && 
b[5932] == 5932 && 
b[5933] == 5933 && 
b[5934] == 5934 && 
b[5935] == 5935 && 
b[5936] == 5936 && 
b[5937] == 5937 && 
b[5938] == 5938 && 
b[5939] == 5939 && 
b[5940] == 5940 && 
b[5941] == 5941 && 
b[5942] == 5942 && 
b[5943] == 5943 && 
b[5944] == 5944 && 
b[5945] == 5945 && 
b[5946] == 5946 && 
b[5947] == 5947 && 
b[5948] == 5948 && 
b[5949] == 5949 && 
b[5950] == 5950 && 
b[5951] == 5951 && 
b[5952] == 5952 && 
b[5953] == 5953 && 
b[5954] == 5954 && 
b[5955] == 5955 && 
b[5956] == 5956 && 
b[5957] == 5957 && 
b[5958] == 5958 && 
b[5959] == 5959 && 
b[5960] == 5960 && 
b[5961] == 5961 && 
b[5962] == 5962 && 
b[5963] == 5963 && 
b[5964] == 5964 && 
b[5965] == 5965 && 
b[5966] == 5966 && 
b[5967] == 5967 && 
b[5968] == 5968 && 
b[5969] == 5969 && 
b[5970] == 5970 && 
b[5971] == 5971 && 
b[5972] == 5972 && 
b[5973] == 5973 && 
b[5974] == 5974 && 
b[5975] == 5975 && 
b[5976] == 5976 && 
b[5977] == 5977 && 
b[5978] == 5978 && 
b[5979] == 5979 && 
b[5980] == 5980 && 
b[5981] == 5981 && 
b[5982] == 5982 && 
b[5983] == 5983 && 
b[5984] == 5984 && 
b[5985] == 5985 && 
b[5986] == 5986 && 
b[5987] == 5987 && 
b[5988] == 5988 && 
b[5989] == 5989 && 
b[5990] == 5990 && 
b[5991] == 5991 && 
b[5992] == 5992 && 
b[5993] == 5993 && 
b[5994] == 5994 && 
b[5995] == 5995 && 
b[5996] == 5996 && 
b[5997] == 5997 && 
b[5998] == 5998 && 
b[5999] == 5999 && 
b[6000] == 6000 && 
b[6001] == 6001 && 
b[6002] == 6002 && 
b[6003] == 6003 && 
b[6004] == 6004 && 
b[6005] == 6005 && 
b[6006] == 6006 && 
b[6007] == 6007 && 
b[6008] == 6008 && 
b[6009] == 6009 && 
b[6010] == 6010 && 
b[6011] == 6011 && 
b[6012] == 6012 && 
b[6013] == 6013 && 
b[6014] == 6014 && 
b[6015] == 6015 && 
b[6016] == 6016 && 
b[6017] == 6017 && 
b[6018] == 6018 && 
b[6019] == 6019 && 
b[6020] == 6020 && 
b[6021] == 6021 && 
b[6022] == 6022 && 
b[6023] == 6023 && 
b[6024] == 6024 && 
b[6025] == 6025 && 
b[6026] == 6026 && 
b[6027] == 6027 && 
b[6028] == 6028 && 
b[6029] == 6029 && 
b[6030] == 6030 && 
b[6031] == 6031 && 
b[6032] == 6032 && 
b[6033] == 6033 && 
b[6034] == 6034 && 
b[6035] == 6035 && 
b[6036] == 6036 && 
b[6037] == 6037 && 
b[6038] == 6038 && 
b[6039] == 6039 && 
b[6040] == 6040 && 
b[6041] == 6041 && 
b[6042] == 6042 && 
b[6043] == 6043 && 
b[6044] == 6044 && 
b[6045] == 6045 && 
b[6046] == 6046 && 
b[6047] == 6047 && 
b[6048] == 6048 && 
b[6049] == 6049 && 
b[6050] == 6050 && 
b[6051] == 6051 && 
b[6052] == 6052 && 
b[6053] == 6053 && 
b[6054] == 6054 && 
b[6055] == 6055 && 
b[6056] == 6056 && 
b[6057] == 6057 && 
b[6058] == 6058 && 
b[6059] == 6059 && 
b[6060] == 6060 && 
b[6061] == 6061 && 
b[6062] == 6062 && 
b[6063] == 6063 && 
b[6064] == 6064 && 
b[6065] == 6065 && 
b[6066] == 6066 && 
b[6067] == 6067 && 
b[6068] == 6068 && 
b[6069] == 6069 && 
b[6070] == 6070 && 
b[6071] == 6071 && 
b[6072] == 6072 && 
b[6073] == 6073 && 
b[6074] == 6074 && 
b[6075] == 6075 && 
b[6076] == 6076 && 
b[6077] == 6077 && 
b[6078] == 6078 && 
b[6079] == 6079 && 
b[6080] == 6080 && 
b[6081] == 6081 && 
b[6082] == 6082 && 
b[6083] == 6083 && 
b[6084] == 6084 && 
b[6085] == 6085 && 
b[6086] == 6086 && 
b[6087] == 6087 && 
b[6088] == 6088 && 
b[6089] == 6089 && 
b[6090] == 6090 && 
b[6091] == 6091 && 
b[6092] == 6092 && 
b[6093] == 6093 && 
b[6094] == 6094 && 
b[6095] == 6095 && 
b[6096] == 6096 && 
b[6097] == 6097 && 
b[6098] == 6098 && 
b[6099] == 6099 && 
b[6100] == 6100 && 
b[6101] == 6101 && 
b[6102] == 6102 && 
b[6103] == 6103 && 
b[6104] == 6104 && 
b[6105] == 6105 && 
b[6106] == 6106 && 
b[6107] == 6107 && 
b[6108] == 6108 && 
b[6109] == 6109 && 
b[6110] == 6110 && 
b[6111] == 6111 && 
b[6112] == 6112 && 
b[6113] == 6113 && 
b[6114] == 6114 && 
b[6115] == 6115 && 
b[6116] == 6116 && 
b[6117] == 6117 && 
b[6118] == 6118 && 
b[6119] == 6119 && 
b[6120] == 6120 && 
b[6121] == 6121 && 
b[6122] == 6122 && 
b[6123] == 6123 && 
b[6124] == 6124 && 
b[6125] == 6125 && 
b[6126] == 6126 && 
b[6127] == 6127 && 
b[6128] == 6128 && 
b[6129] == 6129 && 
b[6130] == 6130 && 
b[6131] == 6131 && 
b[6132] == 6132 && 
b[6133] == 6133 && 
b[6134] == 6134 && 
b[6135] == 6135 && 
b[6136] == 6136 && 
b[6137] == 6137 && 
b[6138] == 6138 && 
b[6139] == 6139 && 
b[6140] == 6140 && 
b[6141] == 6141 && 
b[6142] == 6142 && 
b[6143] == 6143 && 
b[6144] == 6144 && 
b[6145] == 6145 && 
b[6146] == 6146 && 
b[6147] == 6147 && 
b[6148] == 6148 && 
b[6149] == 6149 && 
b[6150] == 6150 && 
b[6151] == 6151 && 
b[6152] == 6152 && 
b[6153] == 6153 && 
b[6154] == 6154 && 
b[6155] == 6155 && 
b[6156] == 6156 && 
b[6157] == 6157 && 
b[6158] == 6158 && 
b[6159] == 6159 && 
b[6160] == 6160 && 
b[6161] == 6161 && 
b[6162] == 6162 && 
b[6163] == 6163 && 
b[6164] == 6164 && 
b[6165] == 6165 && 
b[6166] == 6166 && 
b[6167] == 6167 && 
b[6168] == 6168 && 
b[6169] == 6169 && 
b[6170] == 6170 && 
b[6171] == 6171 && 
b[6172] == 6172 && 
b[6173] == 6173 && 
b[6174] == 6174 && 
b[6175] == 6175 && 
b[6176] == 6176 && 
b[6177] == 6177 && 
b[6178] == 6178 && 
b[6179] == 6179 && 
b[6180] == 6180 && 
b[6181] == 6181 && 
b[6182] == 6182 && 
b[6183] == 6183 && 
b[6184] == 6184 && 
b[6185] == 6185 && 
b[6186] == 6186 && 
b[6187] == 6187 && 
b[6188] == 6188 && 
b[6189] == 6189 && 
b[6190] == 6190 && 
b[6191] == 6191 && 
b[6192] == 6192 && 
b[6193] == 6193 && 
b[6194] == 6194 && 
b[6195] == 6195 && 
b[6196] == 6196 && 
b[6197] == 6197 && 
b[6198] == 6198 && 
b[6199] == 6199 && 
b[6200] == 6200 && 
b[6201] == 6201 && 
b[6202] == 6202 && 
b[6203] == 6203 && 
b[6204] == 6204 && 
b[6205] == 6205 && 
b[6206] == 6206 && 
b[6207] == 6207 && 
b[6208] == 6208 && 
b[6209] == 6209 && 
b[6210] == 6210 && 
b[6211] == 6211 && 
b[6212] == 6212 && 
b[6213] == 6213 && 
b[6214] == 6214 && 
b[6215] == 6215 && 
b[6216] == 6216 && 
b[6217] == 6217 && 
b[6218] == 6218 && 
b[6219] == 6219 && 
b[6220] == 6220 && 
b[6221] == 6221 && 
b[6222] == 6222 && 
b[6223] == 6223 && 
b[6224] == 6224 && 
b[6225] == 6225 && 
b[6226] == 6226 && 
b[6227] == 6227 && 
b[6228] == 6228 && 
b[6229] == 6229 && 
b[6230] == 6230 && 
b[6231] == 6231 && 
b[6232] == 6232 && 
b[6233] == 6233 && 
b[6234] == 6234 && 
b[6235] == 6235 && 
b[6236] == 6236 && 
b[6237] == 6237 && 
b[6238] == 6238 && 
b[6239] == 6239 && 
b[6240] == 6240 && 
b[6241] == 6241 && 
b[6242] == 6242 && 
b[6243] == 6243 && 
b[6244] == 6244 && 
b[6245] == 6245 && 
b[6246] == 6246 && 
b[6247] == 6247 && 
b[6248] == 6248 && 
b[6249] == 6249 && 
b[6250] == 6250 && 
b[6251] == 6251 && 
b[6252] == 6252 && 
b[6253] == 6253 && 
b[6254] == 6254 && 
b[6255] == 6255 && 
b[6256] == 6256 && 
b[6257] == 6257 && 
b[6258] == 6258 && 
b[6259] == 6259 && 
b[6260] == 6260 && 
b[6261] == 6261 && 
b[6262] == 6262 && 
b[6263] == 6263 && 
b[6264] == 6264 && 
b[6265] == 6265 && 
b[6266] == 6266 && 
b[6267] == 6267 && 
b[6268] == 6268 && 
b[6269] == 6269 && 
b[6270] == 6270 && 
b[6271] == 6271 && 
b[6272] == 6272 && 
b[6273] == 6273 && 
b[6274] == 6274 && 
b[6275] == 6275 && 
b[6276] == 6276 && 
b[6277] == 6277 && 
b[6278] == 6278 && 
b[6279] == 6279 && 
b[6280] == 6280 && 
b[6281] == 6281 && 
b[6282] == 6282 && 
b[6283] == 6283 && 
b[6284] == 6284 && 
b[6285] == 6285 && 
b[6286] == 6286 && 
b[6287] == 6287 && 
b[6288] == 6288 && 
b[6289] == 6289 && 
b[6290] == 6290 && 
b[6291] == 6291 && 
b[6292] == 6292 && 
b[6293] == 6293 && 
b[6294] == 6294 && 
b[6295] == 6295 && 
b[6296] == 6296 && 
b[6297] == 6297 && 
b[6298] == 6298 && 
b[6299] == 6299 && 
b[6300] == 6300 && 
b[6301] == 6301 && 
b[6302] == 6302 && 
b[6303] == 6303 && 
b[6304] == 6304 && 
b[6305] == 6305 && 
b[6306] == 6306 && 
b[6307] == 6307 && 
b[6308] == 6308 && 
b[6309] == 6309 && 
b[6310] == 6310 && 
b[6311] == 6311 && 
b[6312] == 6312 && 
b[6313] == 6313 && 
b[6314] == 6314 && 
b[6315] == 6315 && 
b[6316] == 6316 && 
b[6317] == 6317 && 
b[6318] == 6318 && 
b[6319] == 6319 && 
b[6320] == 6320 && 
b[6321] == 6321 && 
b[6322] == 6322 && 
b[6323] == 6323 && 
b[6324] == 6324 && 
b[6325] == 6325 && 
b[6326] == 6326 && 
b[6327] == 6327 && 
b[6328] == 6328 && 
b[6329] == 6329 && 
b[6330] == 6330 && 
b[6331] == 6331 && 
b[6332] == 6332 && 
b[6333] == 6333 && 
b[6334] == 6334 && 
b[6335] == 6335 && 
b[6336] == 6336 && 
b[6337] == 6337 && 
b[6338] == 6338 && 
b[6339] == 6339 && 
b[6340] == 6340 && 
b[6341] == 6341 && 
b[6342] == 6342 && 
b[6343] == 6343 && 
b[6344] == 6344 && 
b[6345] == 6345 && 
b[6346] == 6346 && 
b[6347] == 6347 && 
b[6348] == 6348 && 
b[6349] == 6349 && 
b[6350] == 6350 && 
b[6351] == 6351 && 
b[6352] == 6352 && 
b[6353] == 6353 && 
b[6354] == 6354 && 
b[6355] == 6355 && 
b[6356] == 6356 && 
b[6357] == 6357 && 
b[6358] == 6358 && 
b[6359] == 6359 && 
b[6360] == 6360 && 
b[6361] == 6361 && 
b[6362] == 6362 && 
b[6363] == 6363 && 
b[6364] == 6364 && 
b[6365] == 6365 && 
b[6366] == 6366 && 
b[6367] == 6367 && 
b[6368] == 6368 && 
b[6369] == 6369 && 
b[6370] == 6370 && 
b[6371] == 6371 && 
b[6372] == 6372 && 
b[6373] == 6373 && 
b[6374] == 6374 && 
b[6375] == 6375 && 
b[6376] == 6376 && 
b[6377] == 6377 && 
b[6378] == 6378 && 
b[6379] == 6379 && 
b[6380] == 6380 && 
b[6381] == 6381 && 
b[6382] == 6382 && 
b[6383] == 6383 && 
b[6384] == 6384 && 
b[6385] == 6385 && 
b[6386] == 6386 && 
b[6387] == 6387 && 
b[6388] == 6388 && 
b[6389] == 6389 && 
b[6390] == 6390 && 
b[6391] == 6391 && 
b[6392] == 6392 && 
b[6393] == 6393 && 
b[6394] == 6394 && 
b[6395] == 6395 && 
b[6396] == 6396 && 
b[6397] == 6397 && 
b[6398] == 6398 && 
b[6399] == 6399 && 
b[6400] == 6400 && 
b[6401] == 6401 && 
b[6402] == 6402 && 
b[6403] == 6403 && 
b[6404] == 6404 && 
b[6405] == 6405 && 
b[6406] == 6406 && 
b[6407] == 6407 && 
b[6408] == 6408 && 
b[6409] == 6409 && 
b[6410] == 6410 && 
b[6411] == 6411 && 
b[6412] == 6412 && 
b[6413] == 6413 && 
b[6414] == 6414 && 
b[6415] == 6415 && 
b[6416] == 6416 && 
b[6417] == 6417 && 
b[6418] == 6418 && 
b[6419] == 6419 && 
b[6420] == 6420 && 
b[6421] == 6421 && 
b[6422] == 6422 && 
b[6423] == 6423 && 
b[6424] == 6424 && 
b[6425] == 6425 && 
b[6426] == 6426 && 
b[6427] == 6427 && 
b[6428] == 6428 && 
b[6429] == 6429 && 
b[6430] == 6430 && 
b[6431] == 6431 && 
b[6432] == 6432 && 
b[6433] == 6433 && 
b[6434] == 6434 && 
b[6435] == 6435 && 
b[6436] == 6436 && 
b[6437] == 6437 && 
b[6438] == 6438 && 
b[6439] == 6439 && 
b[6440] == 6440 && 
b[6441] == 6441 && 
b[6442] == 6442 && 
b[6443] == 6443 && 
b[6444] == 6444 && 
b[6445] == 6445 && 
b[6446] == 6446 && 
b[6447] == 6447 && 
b[6448] == 6448 && 
b[6449] == 6449 && 
b[6450] == 6450 && 
b[6451] == 6451 && 
b[6452] == 6452 && 
b[6453] == 6453 && 
b[6454] == 6454 && 
b[6455] == 6455 && 
b[6456] == 6456 && 
b[6457] == 6457 && 
b[6458] == 6458 && 
b[6459] == 6459 && 
b[6460] == 6460 && 
b[6461] == 6461 && 
b[6462] == 6462 && 
b[6463] == 6463 && 
b[6464] == 6464 && 
b[6465] == 6465 && 
b[6466] == 6466 && 
b[6467] == 6467 && 
b[6468] == 6468 && 
b[6469] == 6469 && 
b[6470] == 6470 && 
b[6471] == 6471 && 
b[6472] == 6472 && 
b[6473] == 6473 && 
b[6474] == 6474 && 
b[6475] == 6475 && 
b[6476] == 6476 && 
b[6477] == 6477 && 
b[6478] == 6478 && 
b[6479] == 6479 && 
b[6480] == 6480 && 
b[6481] == 6481 && 
b[6482] == 6482 && 
b[6483] == 6483 && 
b[6484] == 6484 && 
b[6485] == 6485 && 
b[6486] == 6486 && 
b[6487] == 6487 && 
b[6488] == 6488 && 
b[6489] == 6489 && 
b[6490] == 6490 && 
b[6491] == 6491 && 
b[6492] == 6492 && 
b[6493] == 6493 && 
b[6494] == 6494 && 
b[6495] == 6495 && 
b[6496] == 6496 && 
b[6497] == 6497 && 
b[6498] == 6498 && 
b[6499] == 6499 && 
b[6500] == 6500 && 
b[6501] == 6501 && 
b[6502] == 6502 && 
b[6503] == 6503 && 
b[6504] == 6504 && 
b[6505] == 6505 && 
b[6506] == 6506 && 
b[6507] == 6507 && 
b[6508] == 6508 && 
b[6509] == 6509 && 
b[6510] == 6510 && 
b[6511] == 6511 && 
b[6512] == 6512 && 
b[6513] == 6513 && 
b[6514] == 6514 && 
b[6515] == 6515 && 
b[6516] == 6516 && 
b[6517] == 6517 && 
b[6518] == 6518 && 
b[6519] == 6519 && 
b[6520] == 6520 && 
b[6521] == 6521 && 
b[6522] == 6522 && 
b[6523] == 6523 && 
b[6524] == 6524 && 
b[6525] == 6525 && 
b[6526] == 6526 && 
b[6527] == 6527 && 
b[6528] == 6528 && 
b[6529] == 6529 && 
b[6530] == 6530 && 
b[6531] == 6531 && 
b[6532] == 6532 && 
b[6533] == 6533 && 
b[6534] == 6534 && 
b[6535] == 6535 && 
b[6536] == 6536 && 
b[6537] == 6537 && 
b[6538] == 6538 && 
b[6539] == 6539 && 
b[6540] == 6540 && 
b[6541] == 6541 && 
b[6542] == 6542 && 
b[6543] == 6543 && 
b[6544] == 6544 && 
b[6545] == 6545 && 
b[6546] == 6546 && 
b[6547] == 6547 && 
b[6548] == 6548 && 
b[6549] == 6549 && 
b[6550] == 6550 && 
b[6551] == 6551 && 
b[6552] == 6552 && 
b[6553] == 6553 && 
b[6554] == 6554 && 
b[6555] == 6555 && 
b[6556] == 6556 && 
b[6557] == 6557 && 
b[6558] == 6558 && 
b[6559] == 6559 && 
b[6560] == 6560 && 
b[6561] == 6561 && 
b[6562] == 6562 && 
b[6563] == 6563 && 
b[6564] == 6564 && 
b[6565] == 6565 && 
b[6566] == 6566 && 
b[6567] == 6567 && 
b[6568] == 6568 && 
b[6569] == 6569 && 
b[6570] == 6570 && 
b[6571] == 6571 && 
b[6572] == 6572 && 
b[6573] == 6573 && 
b[6574] == 6574 && 
b[6575] == 6575 && 
b[6576] == 6576 && 
b[6577] == 6577 && 
b[6578] == 6578 && 
b[6579] == 6579 && 
b[6580] == 6580 && 
b[6581] == 6581 && 
b[6582] == 6582 && 
b[6583] == 6583 && 
b[6584] == 6584 && 
b[6585] == 6585 && 
b[6586] == 6586 && 
b[6587] == 6587 && 
b[6588] == 6588 && 
b[6589] == 6589 && 
b[6590] == 6590 && 
b[6591] == 6591 && 
b[6592] == 6592 && 
b[6593] == 6593 && 
b[6594] == 6594 && 
b[6595] == 6595 && 
b[6596] == 6596 && 
b[6597] == 6597 && 
b[6598] == 6598 && 
b[6599] == 6599 && 
b[6600] == 6600 && 
b[6601] == 6601 && 
b[6602] == 6602 && 
b[6603] == 6603 && 
b[6604] == 6604 && 
b[6605] == 6605 && 
b[6606] == 6606 && 
b[6607] == 6607 && 
b[6608] == 6608 && 
b[6609] == 6609 && 
b[6610] == 6610 && 
b[6611] == 6611 && 
b[6612] == 6612 && 
b[6613] == 6613 && 
b[6614] == 6614 && 
b[6615] == 6615 && 
b[6616] == 6616 && 
b[6617] == 6617 && 
b[6618] == 6618 && 
b[6619] == 6619 && 
b[6620] == 6620 && 
b[6621] == 6621 && 
b[6622] == 6622 && 
b[6623] == 6623 && 
b[6624] == 6624 && 
b[6625] == 6625 && 
b[6626] == 6626 && 
b[6627] == 6627 && 
b[6628] == 6628 && 
b[6629] == 6629 && 
b[6630] == 6630 && 
b[6631] == 6631 && 
b[6632] == 6632 && 
b[6633] == 6633 && 
b[6634] == 6634 && 
b[6635] == 6635 && 
b[6636] == 6636 && 
b[6637] == 6637 && 
b[6638] == 6638 && 
b[6639] == 6639 && 
b[6640] == 6640 && 
b[6641] == 6641 && 
b[6642] == 6642 && 
b[6643] == 6643 && 
b[6644] == 6644 && 
b[6645] == 6645 && 
b[6646] == 6646 && 
b[6647] == 6647 && 
b[6648] == 6648 && 
b[6649] == 6649 && 
b[6650] == 6650 && 
b[6651] == 6651 && 
b[6652] == 6652 && 
b[6653] == 6653 && 
b[6654] == 6654 && 
b[6655] == 6655 && 
b[6656] == 6656 && 
b[6657] == 6657 && 
b[6658] == 6658 && 
b[6659] == 6659 && 
b[6660] == 6660 && 
b[6661] == 6661 && 
b[6662] == 6662 && 
b[6663] == 6663 && 
b[6664] == 6664 && 
b[6665] == 6665 && 
b[6666] == 6666 && 
b[6667] == 6667 && 
b[6668] == 6668 && 
b[6669] == 6669 && 
b[6670] == 6670 && 
b[6671] == 6671 && 
b[6672] == 6672 && 
b[6673] == 6673 && 
b[6674] == 6674 && 
b[6675] == 6675 && 
b[6676] == 6676 && 
b[6677] == 6677 && 
b[6678] == 6678 && 
b[6679] == 6679 && 
b[6680] == 6680 && 
b[6681] == 6681 && 
b[6682] == 6682 && 
b[6683] == 6683 && 
b[6684] == 6684 && 
b[6685] == 6685 && 
b[6686] == 6686 && 
b[6687] == 6687 && 
b[6688] == 6688 && 
b[6689] == 6689 && 
b[6690] == 6690 && 
b[6691] == 6691 && 
b[6692] == 6692 && 
b[6693] == 6693 && 
b[6694] == 6694 && 
b[6695] == 6695 && 
b[6696] == 6696 && 
b[6697] == 6697 && 
b[6698] == 6698 && 
b[6699] == 6699 && 
b[6700] == 6700 && 
b[6701] == 6701 && 
b[6702] == 6702 && 
b[6703] == 6703 && 
b[6704] == 6704 && 
b[6705] == 6705 && 
b[6706] == 6706 && 
b[6707] == 6707 && 
b[6708] == 6708 && 
b[6709] == 6709 && 
b[6710] == 6710 && 
b[6711] == 6711 && 
b[6712] == 6712 && 
b[6713] == 6713 && 
b[6714] == 6714 && 
b[6715] == 6715 && 
b[6716] == 6716 && 
b[6717] == 6717 && 
b[6718] == 6718 && 
b[6719] == 6719 && 
b[6720] == 6720 && 
b[6721] == 6721 && 
b[6722] == 6722 && 
b[6723] == 6723 && 
b[6724] == 6724 && 
b[6725] == 6725 && 
b[6726] == 6726 && 
b[6727] == 6727 && 
b[6728] == 6728 && 
b[6729] == 6729 && 
b[6730] == 6730 && 
b[6731] == 6731 && 
b[6732] == 6732 && 
b[6733] == 6733 && 
b[6734] == 6734 && 
b[6735] == 6735 && 
b[6736] == 6736 && 
b[6737] == 6737 && 
b[6738] == 6738 && 
b[6739] == 6739 && 
b[6740] == 6740 && 
b[6741] == 6741 && 
b[6742] == 6742 && 
b[6743] == 6743 && 
b[6744] == 6744 && 
b[6745] == 6745 && 
b[6746] == 6746 && 
b[6747] == 6747 && 
b[6748] == 6748 && 
b[6749] == 6749 && 
b[6750] == 6750 && 
b[6751] == 6751 && 
b[6752] == 6752 && 
b[6753] == 6753 && 
b[6754] == 6754 && 
b[6755] == 6755 && 
b[6756] == 6756 && 
b[6757] == 6757 && 
b[6758] == 6758 && 
b[6759] == 6759 && 
b[6760] == 6760 && 
b[6761] == 6761 && 
b[6762] == 6762 && 
b[6763] == 6763 && 
b[6764] == 6764 && 
b[6765] == 6765 && 
b[6766] == 6766 && 
b[6767] == 6767 && 
b[6768] == 6768 && 
b[6769] == 6769 && 
b[6770] == 6770 && 
b[6771] == 6771 && 
b[6772] == 6772 && 
b[6773] == 6773 && 
b[6774] == 6774 && 
b[6775] == 6775 && 
b[6776] == 6776 && 
b[6777] == 6777 && 
b[6778] == 6778 && 
b[6779] == 6779 && 
b[6780] == 6780 && 
b[6781] == 6781 && 
b[6782] == 6782 && 
b[6783] == 6783 && 
b[6784] == 6784 && 
b[6785] == 6785 && 
b[6786] == 6786 && 
b[6787] == 6787 && 
b[6788] == 6788 && 
b[6789] == 6789 && 
b[6790] == 6790 && 
b[6791] == 6791 && 
b[6792] == 6792 && 
b[6793] == 6793 && 
b[6794] == 6794 && 
b[6795] == 6795 && 
b[6796] == 6796 && 
b[6797] == 6797 && 
b[6798] == 6798 && 
b[6799] == 6799 && 
b[6800] == 6800 && 
b[6801] == 6801 && 
b[6802] == 6802 && 
b[6803] == 6803 && 
b[6804] == 6804 && 
b[6805] == 6805 && 
b[6806] == 6806 && 
b[6807] == 6807 && 
b[6808] == 6808 && 
b[6809] == 6809 && 
b[6810] == 6810 && 
b[6811] == 6811 && 
b[6812] == 6812 && 
b[6813] == 6813 && 
b[6814] == 6814 && 
b[6815] == 6815 && 
b[6816] == 6816 && 
b[6817] == 6817 && 
b[6818] == 6818 && 
b[6819] == 6819 && 
b[6820] == 6820 && 
b[6821] == 6821 && 
b[6822] == 6822 && 
b[6823] == 6823 && 
b[6824] == 6824 && 
b[6825] == 6825 && 
b[6826] == 6826 && 
b[6827] == 6827 && 
b[6828] == 6828 && 
b[6829] == 6829 && 
b[6830] == 6830 && 
b[6831] == 6831 && 
b[6832] == 6832 && 
b[6833] == 6833 && 
b[6834] == 6834 && 
b[6835] == 6835 && 
b[6836] == 6836 && 
b[6837] == 6837 && 
b[6838] == 6838 && 
b[6839] == 6839 && 
b[6840] == 6840 && 
b[6841] == 6841 && 
b[6842] == 6842 && 
b[6843] == 6843 && 
b[6844] == 6844 && 
b[6845] == 6845 && 
b[6846] == 6846 && 
b[6847] == 6847 && 
b[6848] == 6848 && 
b[6849] == 6849 && 
b[6850] == 6850 && 
b[6851] == 6851 && 
b[6852] == 6852 && 
b[6853] == 6853 && 
b[6854] == 6854 && 
b[6855] == 6855 && 
b[6856] == 6856 && 
b[6857] == 6857 && 
b[6858] == 6858 && 
b[6859] == 6859 && 
b[6860] == 6860 && 
b[6861] == 6861 && 
b[6862] == 6862 && 
b[6863] == 6863 && 
b[6864] == 6864 && 
b[6865] == 6865 && 
b[6866] == 6866 && 
b[6867] == 6867 && 
b[6868] == 6868 && 
b[6869] == 6869 && 
b[6870] == 6870 && 
b[6871] == 6871 && 
b[6872] == 6872 && 
b[6873] == 6873 && 
b[6874] == 6874 && 
b[6875] == 6875 && 
b[6876] == 6876 && 
b[6877] == 6877 && 
b[6878] == 6878 && 
b[6879] == 6879 && 
b[6880] == 6880 && 
b[6881] == 6881 && 
b[6882] == 6882 && 
b[6883] == 6883 && 
b[6884] == 6884 && 
b[6885] == 6885 && 
b[6886] == 6886 && 
b[6887] == 6887 && 
b[6888] == 6888 && 
b[6889] == 6889 && 
b[6890] == 6890 && 
b[6891] == 6891 && 
b[6892] == 6892 && 
b[6893] == 6893 && 
b[6894] == 6894 && 
b[6895] == 6895 && 
b[6896] == 6896 && 
b[6897] == 6897 && 
b[6898] == 6898 && 
b[6899] == 6899 && 
b[6900] == 6900 && 
b[6901] == 6901 && 
b[6902] == 6902 && 
b[6903] == 6903 && 
b[6904] == 6904 && 
b[6905] == 6905 && 
b[6906] == 6906 && 
b[6907] == 6907 && 
b[6908] == 6908 && 
b[6909] == 6909 && 
b[6910] == 6910 && 
b[6911] == 6911 && 
b[6912] == 6912 && 
b[6913] == 6913 && 
b[6914] == 6914 && 
b[6915] == 6915 && 
b[6916] == 6916 && 
b[6917] == 6917 && 
b[6918] == 6918 && 
b[6919] == 6919 && 
b[6920] == 6920 && 
b[6921] == 6921 && 
b[6922] == 6922 && 
b[6923] == 6923 && 
b[6924] == 6924 && 
b[6925] == 6925 && 
b[6926] == 6926 && 
b[6927] == 6927 && 
b[6928] == 6928 && 
b[6929] == 6929 && 
b[6930] == 6930 && 
b[6931] == 6931 && 
b[6932] == 6932 && 
b[6933] == 6933 && 
b[6934] == 6934 && 
b[6935] == 6935 && 
b[6936] == 6936 && 
b[6937] == 6937 && 
b[6938] == 6938 && 
b[6939] == 6939 && 
b[6940] == 6940 && 
b[6941] == 6941 && 
b[6942] == 6942 && 
b[6943] == 6943 && 
b[6944] == 6944 && 
b[6945] == 6945 && 
b[6946] == 6946 && 
b[6947] == 6947 && 
b[6948] == 6948 && 
b[6949] == 6949 && 
b[6950] == 6950 && 
b[6951] == 6951 && 
b[6952] == 6952 && 
b[6953] == 6953 && 
b[6954] == 6954 && 
b[6955] == 6955 && 
b[6956] == 6956 && 
b[6957] == 6957 && 
b[6958] == 6958 && 
b[6959] == 6959 && 
b[6960] == 6960 && 
b[6961] == 6961 && 
b[6962] == 6962 && 
b[6963] == 6963 && 
b[6964] == 6964 && 
b[6965] == 6965 && 
b[6966] == 6966 && 
b[6967] == 6967 && 
b[6968] == 6968 && 
b[6969] == 6969 && 
b[6970] == 6970 && 
b[6971] == 6971 && 
b[6972] == 6972 && 
b[6973] == 6973 && 
b[6974] == 6974 && 
b[6975] == 6975 && 
b[6976] == 6976 && 
b[6977] == 6977 && 
b[6978] == 6978 && 
b[6979] == 6979 && 
b[6980] == 6980 && 
b[6981] == 6981 && 
b[6982] == 6982 && 
b[6983] == 6983 && 
b[6984] == 6984 && 
b[6985] == 6985 && 
b[6986] == 6986 && 
b[6987] == 6987 && 
b[6988] == 6988 && 
b[6989] == 6989 && 
b[6990] == 6990 && 
b[6991] == 6991 && 
b[6992] == 6992 && 
b[6993] == 6993 && 
b[6994] == 6994 && 
b[6995] == 6995 && 
b[6996] == 6996 && 
b[6997] == 6997 && 
b[6998] == 6998 && 
b[6999] == 6999 && 
b[7000] == 7000 && 
b[7001] == 7001 && 
b[7002] == 7002 && 
b[7003] == 7003 && 
b[7004] == 7004 && 
b[7005] == 7005 && 
b[7006] == 7006 && 
b[7007] == 7007 && 
b[7008] == 7008 && 
b[7009] == 7009 && 
b[7010] == 7010 && 
b[7011] == 7011 && 
b[7012] == 7012 && 
b[7013] == 7013 && 
b[7014] == 7014 && 
b[7015] == 7015 && 
b[7016] == 7016 && 
b[7017] == 7017 && 
b[7018] == 7018 && 
b[7019] == 7019 && 
b[7020] == 7020 && 
b[7021] == 7021 && 
b[7022] == 7022 && 
b[7023] == 7023 && 
b[7024] == 7024 && 
b[7025] == 7025 && 
b[7026] == 7026 && 
b[7027] == 7027 && 
b[7028] == 7028 && 
b[7029] == 7029 && 
b[7030] == 7030 && 
b[7031] == 7031 && 
b[7032] == 7032 && 
b[7033] == 7033 && 
b[7034] == 7034 && 
b[7035] == 7035 && 
b[7036] == 7036 && 
b[7037] == 7037 && 
b[7038] == 7038 && 
b[7039] == 7039 && 
b[7040] == 7040 && 
b[7041] == 7041 && 
b[7042] == 7042 && 
b[7043] == 7043 && 
b[7044] == 7044 && 
b[7045] == 7045 && 
b[7046] == 7046 && 
b[7047] == 7047 && 
b[7048] == 7048 && 
b[7049] == 7049 && 
b[7050] == 7050 && 
b[7051] == 7051 && 
b[7052] == 7052 && 
b[7053] == 7053 && 
b[7054] == 7054 && 
b[7055] == 7055 && 
b[7056] == 7056 && 
b[7057] == 7057 && 
b[7058] == 7058 && 
b[7059] == 7059 && 
b[7060] == 7060 && 
b[7061] == 7061 && 
b[7062] == 7062 && 
b[7063] == 7063 && 
b[7064] == 7064 && 
b[7065] == 7065 && 
b[7066] == 7066 && 
b[7067] == 7067 && 
b[7068] == 7068 && 
b[7069] == 7069 && 
b[7070] == 7070 && 
b[7071] == 7071 && 
b[7072] == 7072 && 
b[7073] == 7073 && 
b[7074] == 7074 && 
b[7075] == 7075 && 
b[7076] == 7076 && 
b[7077] == 7077 && 
b[7078] == 7078 && 
b[7079] == 7079 && 
b[7080] == 7080 && 
b[7081] == 7081 && 
b[7082] == 7082 && 
b[7083] == 7083 && 
b[7084] == 7084 && 
b[7085] == 7085 && 
b[7086] == 7086 && 
b[7087] == 7087 && 
b[7088] == 7088 && 
b[7089] == 7089 && 
b[7090] == 7090 && 
b[7091] == 7091 && 
b[7092] == 7092 && 
b[7093] == 7093 && 
b[7094] == 7094 && 
b[7095] == 7095 && 
b[7096] == 7096 && 
b[7097] == 7097 && 
b[7098] == 7098 && 
b[7099] == 7099 && 
b[7100] == 7100 && 
b[7101] == 7101 && 
b[7102] == 7102 && 
b[7103] == 7103 && 
b[7104] == 7104 && 
b[7105] == 7105 && 
b[7106] == 7106 && 
b[7107] == 7107 && 
b[7108] == 7108 && 
b[7109] == 7109 && 
b[7110] == 7110 && 
b[7111] == 7111 && 
b[7112] == 7112 && 
b[7113] == 7113 && 
b[7114] == 7114 && 
b[7115] == 7115 && 
b[7116] == 7116 && 
b[7117] == 7117 && 
b[7118] == 7118 && 
b[7119] == 7119 && 
b[7120] == 7120 && 
b[7121] == 7121 && 
b[7122] == 7122 && 
b[7123] == 7123 && 
b[7124] == 7124 && 
b[7125] == 7125 && 
b[7126] == 7126 && 
b[7127] == 7127 && 
b[7128] == 7128 && 
b[7129] == 7129 && 
b[7130] == 7130 && 
b[7131] == 7131 && 
b[7132] == 7132 && 
b[7133] == 7133 && 
b[7134] == 7134 && 
b[7135] == 7135 && 
b[7136] == 7136 && 
b[7137] == 7137 && 
b[7138] == 7138 && 
b[7139] == 7139 && 
b[7140] == 7140 && 
b[7141] == 7141 && 
b[7142] == 7142 && 
b[7143] == 7143 && 
b[7144] == 7144 && 
b[7145] == 7145 && 
b[7146] == 7146 && 
b[7147] == 7147 && 
b[7148] == 7148 && 
b[7149] == 7149 && 
b[7150] == 7150 && 
b[7151] == 7151 && 
b[7152] == 7152 && 
b[7153] == 7153 && 
b[7154] == 7154 && 
b[7155] == 7155 && 
b[7156] == 7156 && 
b[7157] == 7157 && 
b[7158] == 7158 && 
b[7159] == 7159 && 
b[7160] == 7160 && 
b[7161] == 7161 && 
b[7162] == 7162 && 
b[7163] == 7163 && 
b[7164] == 7164 && 
b[7165] == 7165 && 
b[7166] == 7166 && 
b[7167] == 7167 && 
b[7168] == 7168 && 
b[7169] == 7169 && 
b[7170] == 7170 && 
b[7171] == 7171 && 
b[7172] == 7172 && 
b[7173] == 7173 && 
b[7174] == 7174 && 
b[7175] == 7175 && 
b[7176] == 7176 && 
b[7177] == 7177 && 
b[7178] == 7178 && 
b[7179] == 7179 && 
b[7180] == 7180 && 
b[7181] == 7181 && 
b[7182] == 7182 && 
b[7183] == 7183 && 
b[7184] == 7184 && 
b[7185] == 7185 && 
b[7186] == 7186 && 
b[7187] == 7187 && 
b[7188] == 7188 && 
b[7189] == 7189 && 
b[7190] == 7190 && 
b[7191] == 7191 && 
b[7192] == 7192 && 
b[7193] == 7193 && 
b[7194] == 7194 && 
b[7195] == 7195 && 
b[7196] == 7196 && 
b[7197] == 7197 && 
b[7198] == 7198 && 
b[7199] == 7199 && 
b[7200] == 7200 && 
b[7201] == 7201 && 
b[7202] == 7202 && 
b[7203] == 7203 && 
b[7204] == 7204 && 
b[7205] == 7205 && 
b[7206] == 7206 && 
b[7207] == 7207 && 
b[7208] == 7208 && 
b[7209] == 7209 && 
b[7210] == 7210 && 
b[7211] == 7211 && 
b[7212] == 7212 && 
b[7213] == 7213 && 
b[7214] == 7214 && 
b[7215] == 7215 && 
b[7216] == 7216 && 
b[7217] == 7217 && 
b[7218] == 7218 && 
b[7219] == 7219 && 
b[7220] == 7220 && 
b[7221] == 7221 && 
b[7222] == 7222 && 
b[7223] == 7223 && 
b[7224] == 7224 && 
b[7225] == 7225 && 
b[7226] == 7226 && 
b[7227] == 7227 && 
b[7228] == 7228 && 
b[7229] == 7229 && 
b[7230] == 7230 && 
b[7231] == 7231 && 
b[7232] == 7232 && 
b[7233] == 7233 && 
b[7234] == 7234 && 
b[7235] == 7235 && 
b[7236] == 7236 && 
b[7237] == 7237 && 
b[7238] == 7238 && 
b[7239] == 7239 && 
b[7240] == 7240 && 
b[7241] == 7241 && 
b[7242] == 7242 && 
b[7243] == 7243 && 
b[7244] == 7244 && 
b[7245] == 7245 && 
b[7246] == 7246 && 
b[7247] == 7247 && 
b[7248] == 7248 && 
b[7249] == 7249 && 
b[7250] == 7250 && 
b[7251] == 7251 && 
b[7252] == 7252 && 
b[7253] == 7253 && 
b[7254] == 7254 && 
b[7255] == 7255 && 
b[7256] == 7256 && 
b[7257] == 7257 && 
b[7258] == 7258 && 
b[7259] == 7259 && 
b[7260] == 7260 && 
b[7261] == 7261 && 
b[7262] == 7262 && 
b[7263] == 7263 && 
b[7264] == 7264 && 
b[7265] == 7265 && 
b[7266] == 7266 && 
b[7267] == 7267 && 
b[7268] == 7268 && 
b[7269] == 7269 && 
b[7270] == 7270 && 
b[7271] == 7271 && 
b[7272] == 7272 && 
b[7273] == 7273 && 
b[7274] == 7274 && 
b[7275] == 7275 && 
b[7276] == 7276 && 
b[7277] == 7277 && 
b[7278] == 7278 && 
b[7279] == 7279 && 
b[7280] == 7280 && 
b[7281] == 7281 && 
b[7282] == 7282 && 
b[7283] == 7283 && 
b[7284] == 7284 && 
b[7285] == 7285 && 
b[7286] == 7286 && 
b[7287] == 7287 && 
b[7288] == 7288 && 
b[7289] == 7289 && 
b[7290] == 7290 && 
b[7291] == 7291 && 
b[7292] == 7292 && 
b[7293] == 7293 && 
b[7294] == 7294 && 
b[7295] == 7295 && 
b[7296] == 7296 && 
b[7297] == 7297 && 
b[7298] == 7298 && 
b[7299] == 7299 && 
b[7300] == 7300 && 
b[7301] == 7301 && 
b[7302] == 7302 && 
b[7303] == 7303 && 
b[7304] == 7304 && 
b[7305] == 7305 && 
b[7306] == 7306 && 
b[7307] == 7307 && 
b[7308] == 7308 && 
b[7309] == 7309 && 
b[7310] == 7310 && 
b[7311] == 7311 && 
b[7312] == 7312 && 
b[7313] == 7313 && 
b[7314] == 7314 && 
b[7315] == 7315 && 
b[7316] == 7316 && 
b[7317] == 7317 && 
b[7318] == 7318 && 
b[7319] == 7319 && 
b[7320] == 7320 && 
b[7321] == 7321 && 
b[7322] == 7322 && 
b[7323] == 7323 && 
b[7324] == 7324 && 
b[7325] == 7325 && 
b[7326] == 7326 && 
b[7327] == 7327 && 
b[7328] == 7328 && 
b[7329] == 7329 && 
b[7330] == 7330 && 
b[7331] == 7331 && 
b[7332] == 7332 && 
b[7333] == 7333 && 
b[7334] == 7334 && 
b[7335] == 7335 && 
b[7336] == 7336 && 
b[7337] == 7337 && 
b[7338] == 7338 && 
b[7339] == 7339 && 
b[7340] == 7340 && 
b[7341] == 7341 && 
b[7342] == 7342 && 
b[7343] == 7343 && 
b[7344] == 7344 && 
b[7345] == 7345 && 
b[7346] == 7346 && 
b[7347] == 7347 && 
b[7348] == 7348 && 
b[7349] == 7349 && 
b[7350] == 7350 && 
b[7351] == 7351 && 
b[7352] == 7352 && 
b[7353] == 7353 && 
b[7354] == 7354 && 
b[7355] == 7355 && 
b[7356] == 7356 && 
b[7357] == 7357 && 
b[7358] == 7358 && 
b[7359] == 7359 && 
b[7360] == 7360 && 
b[7361] == 7361 && 
b[7362] == 7362 && 
b[7363] == 7363 && 
b[7364] == 7364 && 
b[7365] == 7365 && 
b[7366] == 7366 && 
b[7367] == 7367 && 
b[7368] == 7368 && 
b[7369] == 7369 && 
b[7370] == 7370 && 
b[7371] == 7371 && 
b[7372] == 7372 && 
b[7373] == 7373 && 
b[7374] == 7374 && 
b[7375] == 7375 && 
b[7376] == 7376 && 
b[7377] == 7377 && 
b[7378] == 7378 && 
b[7379] == 7379 && 
b[7380] == 7380 && 
b[7381] == 7381 && 
b[7382] == 7382 && 
b[7383] == 7383 && 
b[7384] == 7384 && 
b[7385] == 7385 && 
b[7386] == 7386 && 
b[7387] == 7387 && 
b[7388] == 7388 && 
b[7389] == 7389 && 
b[7390] == 7390 && 
b[7391] == 7391 && 
b[7392] == 7392 && 
b[7393] == 7393 && 
b[7394] == 7394 && 
b[7395] == 7395 && 
b[7396] == 7396 && 
b[7397] == 7397 && 
b[7398] == 7398 && 
b[7399] == 7399 && 
b[7400] == 7400 && 
b[7401] == 7401 && 
b[7402] == 7402 && 
b[7403] == 7403 && 
b[7404] == 7404 && 
b[7405] == 7405 && 
b[7406] == 7406 && 
b[7407] == 7407 && 
b[7408] == 7408 && 
b[7409] == 7409 && 
b[7410] == 7410 && 
b[7411] == 7411 && 
b[7412] == 7412 && 
b[7413] == 7413 && 
b[7414] == 7414 && 
b[7415] == 7415 && 
b[7416] == 7416 && 
b[7417] == 7417 && 
b[7418] == 7418 && 
b[7419] == 7419 && 
b[7420] == 7420 && 
b[7421] == 7421 && 
b[7422] == 7422 && 
b[7423] == 7423 && 
b[7424] == 7424 && 
b[7425] == 7425 && 
b[7426] == 7426 && 
b[7427] == 7427 && 
b[7428] == 7428 && 
b[7429] == 7429 && 
b[7430] == 7430 && 
b[7431] == 7431 && 
b[7432] == 7432 && 
b[7433] == 7433 && 
b[7434] == 7434 && 
b[7435] == 7435 && 
b[7436] == 7436 && 
b[7437] == 7437 && 
b[7438] == 7438 && 
b[7439] == 7439 && 
b[7440] == 7440 && 
b[7441] == 7441 && 
b[7442] == 7442 && 
b[7443] == 7443 && 
b[7444] == 7444 && 
b[7445] == 7445 && 
b[7446] == 7446 && 
b[7447] == 7447 && 
b[7448] == 7448 && 
b[7449] == 7449 && 
b[7450] == 7450 && 
b[7451] == 7451 && 
b[7452] == 7452 && 
b[7453] == 7453 && 
b[7454] == 7454 && 
b[7455] == 7455 && 
b[7456] == 7456 && 
b[7457] == 7457 && 
b[7458] == 7458 && 
b[7459] == 7459 && 
b[7460] == 7460 && 
b[7461] == 7461 && 
b[7462] == 7462 && 
b[7463] == 7463 && 
b[7464] == 7464 && 
b[7465] == 7465 && 
b[7466] == 7466 && 
b[7467] == 7467 && 
b[7468] == 7468 && 
b[7469] == 7469 && 
b[7470] == 7470 && 
b[7471] == 7471 && 
b[7472] == 7472 && 
b[7473] == 7473 && 
b[7474] == 7474 && 
b[7475] == 7475 && 
b[7476] == 7476 && 
b[7477] == 7477 && 
b[7478] == 7478 && 
b[7479] == 7479 && 
b[7480] == 7480 && 
b[7481] == 7481 && 
b[7482] == 7482 && 
b[7483] == 7483 && 
b[7484] == 7484 && 
b[7485] == 7485 && 
b[7486] == 7486 && 
b[7487] == 7487 && 
b[7488] == 7488 && 
b[7489] == 7489 && 
b[7490] == 7490 && 
b[7491] == 7491 && 
b[7492] == 7492 && 
b[7493] == 7493 && 
b[7494] == 7494 && 
b[7495] == 7495 && 
b[7496] == 7496 && 
b[7497] == 7497 && 
b[7498] == 7498 && 
b[7499] == 7499 && 
b[7500] == 7500 && 
b[7501] == 7501 && 
b[7502] == 7502 && 
b[7503] == 7503 && 
b[7504] == 7504 && 
b[7505] == 7505 && 
b[7506] == 7506 && 
b[7507] == 7507 && 
b[7508] == 7508 && 
b[7509] == 7509 && 
b[7510] == 7510 && 
b[7511] == 7511 && 
b[7512] == 7512 && 
b[7513] == 7513 && 
b[7514] == 7514 && 
b[7515] == 7515 && 
b[7516] == 7516 && 
b[7517] == 7517 && 
b[7518] == 7518 && 
b[7519] == 7519 && 
b[7520] == 7520 && 
b[7521] == 7521 && 
b[7522] == 7522 && 
b[7523] == 7523 && 
b[7524] == 7524 && 
b[7525] == 7525 && 
b[7526] == 7526 && 
b[7527] == 7527 && 
b[7528] == 7528 && 
b[7529] == 7529 && 
b[7530] == 7530 && 
b[7531] == 7531 && 
b[7532] == 7532 && 
b[7533] == 7533 && 
b[7534] == 7534 && 
b[7535] == 7535 && 
b[7536] == 7536 && 
b[7537] == 7537 && 
b[7538] == 7538 && 
b[7539] == 7539 && 
b[7540] == 7540 && 
b[7541] == 7541 && 
b[7542] == 7542 && 
b[7543] == 7543 && 
b[7544] == 7544 && 
b[7545] == 7545 && 
b[7546] == 7546 && 
b[7547] == 7547 && 
b[7548] == 7548 && 
b[7549] == 7549 && 
b[7550] == 7550 && 
b[7551] == 7551 && 
b[7552] == 7552 && 
b[7553] == 7553 && 
b[7554] == 7554 && 
b[7555] == 7555 && 
b[7556] == 7556 && 
b[7557] == 7557 && 
b[7558] == 7558 && 
b[7559] == 7559 && 
b[7560] == 7560 && 
b[7561] == 7561 && 
b[7562] == 7562 && 
b[7563] == 7563 && 
b[7564] == 7564 && 
b[7565] == 7565 && 
b[7566] == 7566 && 
b[7567] == 7567 && 
b[7568] == 7568 && 
b[7569] == 7569 && 
b[7570] == 7570 && 
b[7571] == 7571 && 
b[7572] == 7572 && 
b[7573] == 7573 && 
b[7574] == 7574 && 
b[7575] == 7575 && 
b[7576] == 7576 && 
b[7577] == 7577 && 
b[7578] == 7578 && 
b[7579] == 7579 && 
b[7580] == 7580 && 
b[7581] == 7581 && 
b[7582] == 7582 && 
b[7583] == 7583 && 
b[7584] == 7584 && 
b[7585] == 7585 && 
b[7586] == 7586 && 
b[7587] == 7587 && 
b[7588] == 7588 && 
b[7589] == 7589 && 
b[7590] == 7590 && 
b[7591] == 7591 && 
b[7592] == 7592 && 
b[7593] == 7593 && 
b[7594] == 7594 && 
b[7595] == 7595 && 
b[7596] == 7596 && 
b[7597] == 7597 && 
b[7598] == 7598 && 
b[7599] == 7599 && 
b[7600] == 7600 && 
b[7601] == 7601 && 
b[7602] == 7602 && 
b[7603] == 7603 && 
b[7604] == 7604 && 
b[7605] == 7605 && 
b[7606] == 7606 && 
b[7607] == 7607 && 
b[7608] == 7608 && 
b[7609] == 7609 && 
b[7610] == 7610 && 
b[7611] == 7611 && 
b[7612] == 7612 && 
b[7613] == 7613 && 
b[7614] == 7614 && 
b[7615] == 7615 && 
b[7616] == 7616 && 
b[7617] == 7617 && 
b[7618] == 7618 && 
b[7619] == 7619 && 
b[7620] == 7620 && 
b[7621] == 7621 && 
b[7622] == 7622 && 
b[7623] == 7623 && 
b[7624] == 7624 && 
b[7625] == 7625 && 
b[7626] == 7626 && 
b[7627] == 7627 && 
b[7628] == 7628 && 
b[7629] == 7629 && 
b[7630] == 7630 && 
b[7631] == 7631 && 
b[7632] == 7632 && 
b[7633] == 7633 && 
b[7634] == 7634 && 
b[7635] == 7635 && 
b[7636] == 7636 && 
b[7637] == 7637 && 
b[7638] == 7638 && 
b[7639] == 7639 && 
b[7640] == 7640 && 
b[7641] == 7641 && 
b[7642] == 7642 && 
b[7643] == 7643 && 
b[7644] == 7644 && 
b[7645] == 7645 && 
b[7646] == 7646 && 
b[7647] == 7647 && 
b[7648] == 7648 && 
b[7649] == 7649 && 
b[7650] == 7650 && 
b[7651] == 7651 && 
b[7652] == 7652 && 
b[7653] == 7653 && 
b[7654] == 7654 && 
b[7655] == 7655 && 
b[7656] == 7656 && 
b[7657] == 7657 && 
b[7658] == 7658 && 
b[7659] == 7659 && 
b[7660] == 7660 && 
b[7661] == 7661 && 
b[7662] == 7662 && 
b[7663] == 7663 && 
b[7664] == 7664 && 
b[7665] == 7665 && 
b[7666] == 7666 && 
b[7667] == 7667 && 
b[7668] == 7668 && 
b[7669] == 7669 && 
b[7670] == 7670 && 
b[7671] == 7671 && 
b[7672] == 7672 && 
b[7673] == 7673 && 
b[7674] == 7674 && 
b[7675] == 7675 && 
b[7676] == 7676 && 
b[7677] == 7677 && 
b[7678] == 7678 && 
b[7679] == 7679 && 
b[7680] == 7680 && 
b[7681] == 7681 && 
b[7682] == 7682 && 
b[7683] == 7683 && 
b[7684] == 7684 && 
b[7685] == 7685 && 
b[7686] == 7686 && 
b[7687] == 7687 && 
b[7688] == 7688 && 
b[7689] == 7689 && 
b[7690] == 7690 && 
b[7691] == 7691 && 
b[7692] == 7692 && 
b[7693] == 7693 && 
b[7694] == 7694 && 
b[7695] == 7695 && 
b[7696] == 7696 && 
b[7697] == 7697 && 
b[7698] == 7698 && 
b[7699] == 7699 && 
b[7700] == 7700 && 
b[7701] == 7701 && 
b[7702] == 7702 && 
b[7703] == 7703 && 
b[7704] == 7704 && 
b[7705] == 7705 && 
b[7706] == 7706 && 
b[7707] == 7707 && 
b[7708] == 7708 && 
b[7709] == 7709 && 
b[7710] == 7710 && 
b[7711] == 7711 && 
b[7712] == 7712 && 
b[7713] == 7713 && 
b[7714] == 7714 && 
b[7715] == 7715 && 
b[7716] == 7716 && 
b[7717] == 7717 && 
b[7718] == 7718 && 
b[7719] == 7719 && 
b[7720] == 7720 && 
b[7721] == 7721 && 
b[7722] == 7722 && 
b[7723] == 7723 && 
b[7724] == 7724 && 
b[7725] == 7725 && 
b[7726] == 7726 && 
b[7727] == 7727 && 
b[7728] == 7728 && 
b[7729] == 7729 && 
b[7730] == 7730 && 
b[7731] == 7731 && 
b[7732] == 7732 && 
b[7733] == 7733 && 
b[7734] == 7734 && 
b[7735] == 7735 && 
b[7736] == 7736 && 
b[7737] == 7737 && 
b[7738] == 7738 && 
b[7739] == 7739 && 
b[7740] == 7740 && 
b[7741] == 7741 && 
b[7742] == 7742 && 
b[7743] == 7743 && 
b[7744] == 7744 && 
b[7745] == 7745 && 
b[7746] == 7746 && 
b[7747] == 7747 && 
b[7748] == 7748 && 
b[7749] == 7749 && 
b[7750] == 7750 && 
b[7751] == 7751 && 
b[7752] == 7752 && 
b[7753] == 7753 && 
b[7754] == 7754 && 
b[7755] == 7755 && 
b[7756] == 7756 && 
b[7757] == 7757 && 
b[7758] == 7758 && 
b[7759] == 7759 && 
b[7760] == 7760 && 
b[7761] == 7761 && 
b[7762] == 7762 && 
b[7763] == 7763 && 
b[7764] == 7764 && 
b[7765] == 7765 && 
b[7766] == 7766 && 
b[7767] == 7767 && 
b[7768] == 7768 && 
b[7769] == 7769 && 
b[7770] == 7770 && 
b[7771] == 7771 && 
b[7772] == 7772 && 
b[7773] == 7773 && 
b[7774] == 7774 && 
b[7775] == 7775 && 
b[7776] == 7776 && 
b[7777] == 7777 && 
b[7778] == 7778 && 
b[7779] == 7779 && 
b[7780] == 7780 && 
b[7781] == 7781 && 
b[7782] == 7782 && 
b[7783] == 7783 && 
b[7784] == 7784 && 
b[7785] == 7785 && 
b[7786] == 7786 && 
b[7787] == 7787 && 
b[7788] == 7788 && 
b[7789] == 7789 && 
b[7790] == 7790 && 
b[7791] == 7791 && 
b[7792] == 7792 && 
b[7793] == 7793 && 
b[7794] == 7794 && 
b[7795] == 7795 && 
b[7796] == 7796 && 
b[7797] == 7797 && 
b[7798] == 7798 && 
b[7799] == 7799 && 
b[7800] == 7800 && 
b[7801] == 7801 && 
b[7802] == 7802 && 
b[7803] == 7803 && 
b[7804] == 7804 && 
b[7805] == 7805 && 
b[7806] == 7806 && 
b[7807] == 7807 && 
b[7808] == 7808 && 
b[7809] == 7809 && 
b[7810] == 7810 && 
b[7811] == 7811 && 
b[7812] == 7812 && 
b[7813] == 7813 && 
b[7814] == 7814 && 
b[7815] == 7815 && 
b[7816] == 7816 && 
b[7817] == 7817 && 
b[7818] == 7818 && 
b[7819] == 7819 && 
b[7820] == 7820 && 
b[7821] == 7821 && 
b[7822] == 7822 && 
b[7823] == 7823 && 
b[7824] == 7824 && 
b[7825] == 7825 && 
b[7826] == 7826 && 
b[7827] == 7827 && 
b[7828] == 7828 && 
b[7829] == 7829 && 
b[7830] == 7830 && 
b[7831] == 7831 && 
b[7832] == 7832 && 
b[7833] == 7833 && 
b[7834] == 7834 && 
b[7835] == 7835 && 
b[7836] == 7836 && 
b[7837] == 7837 && 
b[7838] == 7838 && 
b[7839] == 7839 && 
b[7840] == 7840 && 
b[7841] == 7841 && 
b[7842] == 7842 && 
b[7843] == 7843 && 
b[7844] == 7844 && 
b[7845] == 7845 && 
b[7846] == 7846 && 
b[7847] == 7847 && 
b[7848] == 7848 && 
b[7849] == 7849 && 
b[7850] == 7850 && 
b[7851] == 7851 && 
b[7852] == 7852 && 
b[7853] == 7853 && 
b[7854] == 7854 && 
b[7855] == 7855 && 
b[7856] == 7856 && 
b[7857] == 7857 && 
b[7858] == 7858 && 
b[7859] == 7859 && 
b[7860] == 7860 && 
b[7861] == 7861 && 
b[7862] == 7862 && 
b[7863] == 7863 && 
b[7864] == 7864 && 
b[7865] == 7865 && 
b[7866] == 7866 && 
b[7867] == 7867 && 
b[7868] == 7868 && 
b[7869] == 7869 && 
b[7870] == 7870 && 
b[7871] == 7871 && 
b[7872] == 7872 && 
b[7873] == 7873 && 
b[7874] == 7874 && 
b[7875] == 7875 && 
b[7876] == 7876 && 
b[7877] == 7877 && 
b[7878] == 7878 && 
b[7879] == 7879 && 
b[7880] == 7880 && 
b[7881] == 7881 && 
b[7882] == 7882 && 
b[7883] == 7883 && 
b[7884] == 7884 && 
b[7885] == 7885 && 
b[7886] == 7886 && 
b[7887] == 7887 && 
b[7888] == 7888 && 
b[7889] == 7889 && 
b[7890] == 7890 && 
b[7891] == 7891 && 
b[7892] == 7892 && 
b[7893] == 7893 && 
b[7894] == 7894 && 
b[7895] == 7895 && 
b[7896] == 7896 && 
b[7897] == 7897 && 
b[7898] == 7898 && 
b[7899] == 7899 && 
b[7900] == 7900 && 
b[7901] == 7901 && 
b[7902] == 7902 && 
b[7903] == 7903 && 
b[7904] == 7904 && 
b[7905] == 7905 && 
b[7906] == 7906 && 
b[7907] == 7907 && 
b[7908] == 7908 && 
b[7909] == 7909 && 
b[7910] == 7910 && 
b[7911] == 7911 && 
b[7912] == 7912 && 
b[7913] == 7913 && 
b[7914] == 7914 && 
b[7915] == 7915 && 
b[7916] == 7916 && 
b[7917] == 7917 && 
b[7918] == 7918 && 
b[7919] == 7919 && 
b[7920] == 7920 && 
b[7921] == 7921 && 
b[7922] == 7922 && 
b[7923] == 7923 && 
b[7924] == 7924 && 
b[7925] == 7925 && 
b[7926] == 7926 && 
b[7927] == 7927 && 
b[7928] == 7928 && 
b[7929] == 7929 && 
b[7930] == 7930 && 
b[7931] == 7931 && 
b[7932] == 7932 && 
b[7933] == 7933 && 
b[7934] == 7934 && 
b[7935] == 7935 && 
b[7936] == 7936 && 
b[7937] == 7937 && 
b[7938] == 7938 && 
b[7939] == 7939 && 
b[7940] == 7940 && 
b[7941] == 7941 && 
b[7942] == 7942 && 
b[7943] == 7943 && 
b[7944] == 7944 && 
b[7945] == 7945 && 
b[7946] == 7946 && 
b[7947] == 7947 && 
b[7948] == 7948 && 
b[7949] == 7949 && 
b[7950] == 7950 && 
b[7951] == 7951 && 
b[7952] == 7952 && 
b[7953] == 7953 && 
b[7954] == 7954 && 
b[7955] == 7955 && 
b[7956] == 7956 && 
b[7957] == 7957 && 
b[7958] == 7958 && 
b[7959] == 7959 && 
b[7960] == 7960 && 
b[7961] == 7961 && 
b[7962] == 7962 && 
b[7963] == 7963 && 
b[7964] == 7964 && 
b[7965] == 7965 && 
b[7966] == 7966 && 
b[7967] == 7967 && 
b[7968] == 7968 && 
b[7969] == 7969 && 
b[7970] == 7970 && 
b[7971] == 7971 && 
b[7972] == 7972 && 
b[7973] == 7973 && 
b[7974] == 7974 && 
b[7975] == 7975 && 
b[7976] == 7976 && 
b[7977] == 7977 && 
b[7978] == 7978 && 
b[7979] == 7979 && 
b[7980] == 7980 && 
b[7981] == 7981 && 
b[7982] == 7982 && 
b[7983] == 7983 && 
b[7984] == 7984 && 
b[7985] == 7985 && 
b[7986] == 7986 && 
b[7987] == 7987 && 
b[7988] == 7988 && 
b[7989] == 7989 && 
b[7990] == 7990 && 
b[7991] == 7991 && 
b[7992] == 7992 && 
b[7993] == 7993 && 
b[7994] == 7994 && 
b[7995] == 7995 && 
b[7996] == 7996 && 
b[7997] == 7997 && 
b[7998] == 7998 && 
b[7999] == 7999 && 
b[8000] == 8000 && 
b[8001] == 8001 && 
b[8002] == 8002 && 
b[8003] == 8003 && 
b[8004] == 8004 && 
b[8005] == 8005 && 
b[8006] == 8006 && 
b[8007] == 8007 && 
b[8008] == 8008 && 
b[8009] == 8009 && 
b[8010] == 8010 && 
b[8011] == 8011 && 
b[8012] == 8012 && 
b[8013] == 8013 && 
b[8014] == 8014 && 
b[8015] == 8015 && 
b[8016] == 8016 && 
b[8017] == 8017 && 
b[8018] == 8018 && 
b[8019] == 8019 && 
b[8020] == 8020 && 
b[8021] == 8021 && 
b[8022] == 8022 && 
b[8023] == 8023 && 
b[8024] == 8024 && 
b[8025] == 8025 && 
b[8026] == 8026 && 
b[8027] == 8027 && 
b[8028] == 8028 && 
b[8029] == 8029 && 
b[8030] == 8030 && 
b[8031] == 8031 && 
b[8032] == 8032 && 
b[8033] == 8033 && 
b[8034] == 8034 && 
b[8035] == 8035 && 
b[8036] == 8036 && 
b[8037] == 8037 && 
b[8038] == 8038 && 
b[8039] == 8039 && 
b[8040] == 8040 && 
b[8041] == 8041 && 
b[8042] == 8042 && 
b[8043] == 8043 && 
b[8044] == 8044 && 
b[8045] == 8045 && 
b[8046] == 8046 && 
b[8047] == 8047 && 
b[8048] == 8048 && 
b[8049] == 8049 && 
b[8050] == 8050 && 
b[8051] == 8051 && 
b[8052] == 8052 && 
b[8053] == 8053 && 
b[8054] == 8054 && 
b[8055] == 8055 && 
b[8056] == 8056 && 
b[8057] == 8057 && 
b[8058] == 8058 && 
b[8059] == 8059 && 
b[8060] == 8060 && 
b[8061] == 8061 && 
b[8062] == 8062 && 
b[8063] == 8063 && 
b[8064] == 8064 && 
b[8065] == 8065 && 
b[8066] == 8066 && 
b[8067] == 8067 && 
b[8068] == 8068 && 
b[8069] == 8069 && 
b[8070] == 8070 && 
b[8071] == 8071 && 
b[8072] == 8072 && 
b[8073] == 8073 && 
b[8074] == 8074 && 
b[8075] == 8075 && 
b[8076] == 8076 && 
b[8077] == 8077 && 
b[8078] == 8078 && 
b[8079] == 8079 && 
b[8080] == 8080 && 
b[8081] == 8081 && 
b[8082] == 8082 && 
b[8083] == 8083 && 
b[8084] == 8084 && 
b[8085] == 8085 && 
b[8086] == 8086 && 
b[8087] == 8087 && 
b[8088] == 8088 && 
b[8089] == 8089 && 
b[8090] == 8090 && 
b[8091] == 8091 && 
b[8092] == 8092 && 
b[8093] == 8093 && 
b[8094] == 8094 && 
b[8095] == 8095 && 
b[8096] == 8096 && 
b[8097] == 8097 && 
b[8098] == 8098 && 
b[8099] == 8099 && 
b[8100] == 8100 && 
b[8101] == 8101 && 
b[8102] == 8102 && 
b[8103] == 8103 && 
b[8104] == 8104 && 
b[8105] == 8105 && 
b[8106] == 8106 && 
b[8107] == 8107 && 
b[8108] == 8108 && 
b[8109] == 8109 && 
b[8110] == 8110 && 
b[8111] == 8111 && 
b[8112] == 8112 && 
b[8113] == 8113 && 
b[8114] == 8114 && 
b[8115] == 8115 && 
b[8116] == 8116 && 
b[8117] == 8117 && 
b[8118] == 8118 && 
b[8119] == 8119 && 
b[8120] == 8120 && 
b[8121] == 8121 && 
b[8122] == 8122 && 
b[8123] == 8123 && 
b[8124] == 8124 && 
b[8125] == 8125 && 
b[8126] == 8126 && 
b[8127] == 8127 && 
b[8128] == 8128 && 
b[8129] == 8129 && 
b[8130] == 8130 && 
b[8131] == 8131 && 
b[8132] == 8132 && 
b[8133] == 8133 && 
b[8134] == 8134 && 
b[8135] == 8135 && 
b[8136] == 8136 && 
b[8137] == 8137 && 
b[8138] == 8138 && 
b[8139] == 8139 && 
b[8140] == 8140 && 
b[8141] == 8141 && 
b[8142] == 8142 && 
b[8143] == 8143 && 
b[8144] == 8144 && 
b[8145] == 8145 && 
b[8146] == 8146 && 
b[8147] == 8147 && 
b[8148] == 8148 && 
b[8149] == 8149 && 
b[8150] == 8150 && 
b[8151] == 8151 && 
b[8152] == 8152 && 
b[8153] == 8153 && 
b[8154] == 8154 && 
b[8155] == 8155 && 
b[8156] == 8156 && 
b[8157] == 8157 && 
b[8158] == 8158 && 
b[8159] == 8159 && 
b[8160] == 8160 && 
b[8161] == 8161 && 
b[8162] == 8162 && 
b[8163] == 8163 && 
b[8164] == 8164 && 
b[8165] == 8165 && 
b[8166] == 8166 && 
b[8167] == 8167 && 
b[8168] == 8168 && 
b[8169] == 8169 && 
b[8170] == 8170 && 
b[8171] == 8171 && 
b[8172] == 8172 && 
b[8173] == 8173 && 
b[8174] == 8174 && 
b[8175] == 8175 && 
b[8176] == 8176 && 
b[8177] == 8177 && 
b[8178] == 8178 && 
b[8179] == 8179 && 
b[8180] == 8180 && 
b[8181] == 8181 && 
b[8182] == 8182 && 
b[8183] == 8183 && 
b[8184] == 8184 && 
b[8185] == 8185 && 
b[8186] == 8186 && 
b[8187] == 8187 && 
b[8188] == 8188 && 
b[8189] == 8189 && 
b[8190] == 8190 && 
b[8191] == 8191 && 
b[8192] == 8192 && 
b[8193] == 8193 && 
b[8194] == 8194 && 
b[8195] == 8195 && 
b[8196] == 8196 && 
b[8197] == 8197 && 
b[8198] == 8198 && 
b[8199] == 8199 && 
b[8200] == 8200 && 
b[8201] == 8201 && 
b[8202] == 8202 && 
b[8203] == 8203 && 
b[8204] == 8204 && 
b[8205] == 8205 && 
b[8206] == 8206 && 
b[8207] == 8207 && 
b[8208] == 8208 && 
b[8209] == 8209 && 
b[8210] == 8210 && 
b[8211] == 8211 && 
b[8212] == 8212 && 
b[8213] == 8213 && 
b[8214] == 8214 && 
b[8215] == 8215 && 
b[8216] == 8216 && 
b[8217] == 8217 && 
b[8218] == 8218 && 
b[8219] == 8219 && 
b[8220] == 8220 && 
b[8221] == 8221 && 
b[8222] == 8222 && 
b[8223] == 8223 && 
b[8224] == 8224 && 
b[8225] == 8225 && 
b[8226] == 8226 && 
b[8227] == 8227 && 
b[8228] == 8228 && 
b[8229] == 8229 && 
b[8230] == 8230 && 
b[8231] == 8231 && 
b[8232] == 8232 && 
b[8233] == 8233 && 
b[8234] == 8234 && 
b[8235] == 8235 && 
b[8236] == 8236 && 
b[8237] == 8237 && 
b[8238] == 8238 && 
b[8239] == 8239 && 
b[8240] == 8240 && 
b[8241] == 8241 && 
b[8242] == 8242 && 
b[8243] == 8243 && 
b[8244] == 8244 && 
b[8245] == 8245 && 
b[8246] == 8246 && 
b[8247] == 8247 && 
b[8248] == 8248 && 
b[8249] == 8249 && 
b[8250] == 8250 && 
b[8251] == 8251 && 
b[8252] == 8252 && 
b[8253] == 8253 && 
b[8254] == 8254 && 
b[8255] == 8255 && 
b[8256] == 8256 && 
b[8257] == 8257 && 
b[8258] == 8258 && 
b[8259] == 8259 && 
b[8260] == 8260 && 
b[8261] == 8261 && 
b[8262] == 8262 && 
b[8263] == 8263 && 
b[8264] == 8264 && 
b[8265] == 8265 && 
b[8266] == 8266 && 
b[8267] == 8267 && 
b[8268] == 8268 && 
b[8269] == 8269 && 
b[8270] == 8270 && 
b[8271] == 8271 && 
b[8272] == 8272 && 
b[8273] == 8273 && 
b[8274] == 8274 && 
b[8275] == 8275 && 
b[8276] == 8276 && 
b[8277] == 8277 && 
b[8278] == 8278 && 
b[8279] == 8279 && 
b[8280] == 8280 && 
b[8281] == 8281 && 
b[8282] == 8282 && 
b[8283] == 8283 && 
b[8284] == 8284 && 
b[8285] == 8285 && 
b[8286] == 8286 && 
b[8287] == 8287 && 
b[8288] == 8288 && 
b[8289] == 8289 && 
b[8290] == 8290 && 
b[8291] == 8291 && 
b[8292] == 8292 && 
b[8293] == 8293 && 
b[8294] == 8294 && 
b[8295] == 8295 && 
b[8296] == 8296 && 
b[8297] == 8297 && 
b[8298] == 8298 && 
b[8299] == 8299 && 
b[8300] == 8300 && 
b[8301] == 8301 && 
b[8302] == 8302 && 
b[8303] == 8303 && 
b[8304] == 8304 && 
b[8305] == 8305 && 
b[8306] == 8306 && 
b[8307] == 8307 && 
b[8308] == 8308 && 
b[8309] == 8309 && 
b[8310] == 8310 && 
b[8311] == 8311 && 
b[8312] == 8312 && 
b[8313] == 8313 && 
b[8314] == 8314 && 
b[8315] == 8315 && 
b[8316] == 8316 && 
b[8317] == 8317 && 
b[8318] == 8318 && 
b[8319] == 8319 && 
b[8320] == 8320 && 
b[8321] == 8321 && 
b[8322] == 8322 && 
b[8323] == 8323 && 
b[8324] == 8324 && 
b[8325] == 8325 && 
b[8326] == 8326 && 
b[8327] == 8327 && 
b[8328] == 8328 && 
b[8329] == 8329 && 
b[8330] == 8330 && 
b[8331] == 8331 && 
b[8332] == 8332 && 
b[8333] == 8333 && 
b[8334] == 8334 && 
b[8335] == 8335 && 
b[8336] == 8336 && 
b[8337] == 8337 && 
b[8338] == 8338 && 
b[8339] == 8339 && 
b[8340] == 8340 && 
b[8341] == 8341 && 
b[8342] == 8342 && 
b[8343] == 8343 && 
b[8344] == 8344 && 
b[8345] == 8345 && 
b[8346] == 8346 && 
b[8347] == 8347 && 
b[8348] == 8348 && 
b[8349] == 8349 && 
b[8350] == 8350 && 
b[8351] == 8351 && 
b[8352] == 8352 && 
b[8353] == 8353 && 
b[8354] == 8354 && 
b[8355] == 8355 && 
b[8356] == 8356 && 
b[8357] == 8357 && 
b[8358] == 8358 && 
b[8359] == 8359 && 
b[8360] == 8360 && 
b[8361] == 8361 && 
b[8362] == 8362 && 
b[8363] == 8363 && 
b[8364] == 8364 && 
b[8365] == 8365 && 
b[8366] == 8366 && 
b[8367] == 8367 && 
b[8368] == 8368 && 
b[8369] == 8369 && 
b[8370] == 8370 && 
b[8371] == 8371 && 
b[8372] == 8372 && 
b[8373] == 8373 && 
b[8374] == 8374 && 
b[8375] == 8375 && 
b[8376] == 8376 && 
b[8377] == 8377 && 
b[8378] == 8378 && 
b[8379] == 8379 && 
b[8380] == 8380 && 
b[8381] == 8381 && 
b[8382] == 8382 && 
b[8383] == 8383 && 
b[8384] == 8384 && 
b[8385] == 8385 && 
b[8386] == 8386 && 
b[8387] == 8387 && 
b[8388] == 8388 && 
b[8389] == 8389 && 
b[8390] == 8390 && 
b[8391] == 8391 && 
b[8392] == 8392 && 
b[8393] == 8393 && 
b[8394] == 8394 && 
b[8395] == 8395 && 
b[8396] == 8396 && 
b[8397] == 8397 && 
b[8398] == 8398 && 
b[8399] == 8399 && 
b[8400] == 8400 && 
b[8401] == 8401 && 
b[8402] == 8402 && 
b[8403] == 8403 && 
b[8404] == 8404 && 
b[8405] == 8405 && 
b[8406] == 8406 && 
b[8407] == 8407 && 
b[8408] == 8408 && 
b[8409] == 8409 && 
b[8410] == 8410 && 
b[8411] == 8411 && 
b[8412] == 8412 && 
b[8413] == 8413 && 
b[8414] == 8414 && 
b[8415] == 8415 && 
b[8416] == 8416 && 
b[8417] == 8417 && 
b[8418] == 8418 && 
b[8419] == 8419 && 
b[8420] == 8420 && 
b[8421] == 8421 && 
b[8422] == 8422 && 
b[8423] == 8423 && 
b[8424] == 8424 && 
b[8425] == 8425 && 
b[8426] == 8426 && 
b[8427] == 8427 && 
b[8428] == 8428 && 
b[8429] == 8429 && 
b[8430] == 8430 && 
b[8431] == 8431 && 
b[8432] == 8432 && 
b[8433] == 8433 && 
b[8434] == 8434 && 
b[8435] == 8435 && 
b[8436] == 8436 && 
b[8437] == 8437 && 
b[8438] == 8438 && 
b[8439] == 8439 && 
b[8440] == 8440 && 
b[8441] == 8441 && 
b[8442] == 8442 && 
b[8443] == 8443 && 
b[8444] == 8444 && 
b[8445] == 8445 && 
b[8446] == 8446 && 
b[8447] == 8447 && 
b[8448] == 8448 && 
b[8449] == 8449 && 
b[8450] == 8450 && 
b[8451] == 8451 && 
b[8452] == 8452 && 
b[8453] == 8453 && 
b[8454] == 8454 && 
b[8455] == 8455 && 
b[8456] == 8456 && 
b[8457] == 8457 && 
b[8458] == 8458 && 
b[8459] == 8459 && 
b[8460] == 8460 && 
b[8461] == 8461 && 
b[8462] == 8462 && 
b[8463] == 8463 && 
b[8464] == 8464 && 
b[8465] == 8465 && 
b[8466] == 8466 && 
b[8467] == 8467 && 
b[8468] == 8468 && 
b[8469] == 8469 && 
b[8470] == 8470 && 
b[8471] == 8471 && 
b[8472] == 8472 && 
b[8473] == 8473 && 
b[8474] == 8474 && 
b[8475] == 8475 && 
b[8476] == 8476 && 
b[8477] == 8477 && 
b[8478] == 8478 && 
b[8479] == 8479 && 
b[8480] == 8480 && 
b[8481] == 8481 && 
b[8482] == 8482 && 
b[8483] == 8483 && 
b[8484] == 8484 && 
b[8485] == 8485 && 
b[8486] == 8486 && 
b[8487] == 8487 && 
b[8488] == 8488 && 
b[8489] == 8489 && 
b[8490] == 8490 && 
b[8491] == 8491 && 
b[8492] == 8492 && 
b[8493] == 8493 && 
b[8494] == 8494 && 
b[8495] == 8495 && 
b[8496] == 8496 && 
b[8497] == 8497 && 
b[8498] == 8498 && 
b[8499] == 8499 && 
b[8500] == 8500 && 
b[8501] == 8501 && 
b[8502] == 8502 && 
b[8503] == 8503 && 
b[8504] == 8504 && 
b[8505] == 8505 && 
b[8506] == 8506 && 
b[8507] == 8507 && 
b[8508] == 8508 && 
b[8509] == 8509 && 
b[8510] == 8510 && 
b[8511] == 8511 && 
b[8512] == 8512 && 
b[8513] == 8513 && 
b[8514] == 8514 && 
b[8515] == 8515 && 
b[8516] == 8516 && 
b[8517] == 8517 && 
b[8518] == 8518 && 
b[8519] == 8519 && 
b[8520] == 8520 && 
b[8521] == 8521 && 
b[8522] == 8522 && 
b[8523] == 8523 && 
b[8524] == 8524 && 
b[8525] == 8525 && 
b[8526] == 8526 && 
b[8527] == 8527 && 
b[8528] == 8528 && 
b[8529] == 8529 && 
b[8530] == 8530 && 
b[8531] == 8531 && 
b[8532] == 8532 && 
b[8533] == 8533 && 
b[8534] == 8534 && 
b[8535] == 8535 && 
b[8536] == 8536 && 
b[8537] == 8537 && 
b[8538] == 8538 && 
b[8539] == 8539 && 
b[8540] == 8540 && 
b[8541] == 8541 && 
b[8542] == 8542 && 
b[8543] == 8543 && 
b[8544] == 8544 && 
b[8545] == 8545 && 
b[8546] == 8546 && 
b[8547] == 8547 && 
b[8548] == 8548 && 
b[8549] == 8549 && 
b[8550] == 8550 && 
b[8551] == 8551 && 
b[8552] == 8552 && 
b[8553] == 8553 && 
b[8554] == 8554 && 
b[8555] == 8555 && 
b[8556] == 8556 && 
b[8557] == 8557 && 
b[8558] == 8558 && 
b[8559] == 8559 && 
b[8560] == 8560 && 
b[8561] == 8561 && 
b[8562] == 8562 && 
b[8563] == 8563 && 
b[8564] == 8564 && 
b[8565] == 8565 && 
b[8566] == 8566 && 
b[8567] == 8567 && 
b[8568] == 8568 && 
b[8569] == 8569 && 
b[8570] == 8570 && 
b[8571] == 8571 && 
b[8572] == 8572 && 
b[8573] == 8573 && 
b[8574] == 8574 && 
b[8575] == 8575 && 
b[8576] == 8576 && 
b[8577] == 8577 && 
b[8578] == 8578 && 
b[8579] == 8579 && 
b[8580] == 8580 && 
b[8581] == 8581 && 
b[8582] == 8582 && 
b[8583] == 8583 && 
b[8584] == 8584 && 
b[8585] == 8585 && 
b[8586] == 8586 && 
b[8587] == 8587 && 
b[8588] == 8588 && 
b[8589] == 8589 && 
b[8590] == 8590 && 
b[8591] == 8591 && 
b[8592] == 8592 && 
b[8593] == 8593 && 
b[8594] == 8594 && 
b[8595] == 8595 && 
b[8596] == 8596 && 
b[8597] == 8597 && 
b[8598] == 8598 && 
b[8599] == 8599 && 
b[8600] == 8600 && 
b[8601] == 8601 && 
b[8602] == 8602 && 
b[8603] == 8603 && 
b[8604] == 8604 && 
b[8605] == 8605 && 
b[8606] == 8606 && 
b[8607] == 8607 && 
b[8608] == 8608 && 
b[8609] == 8609 && 
b[8610] == 8610 && 
b[8611] == 8611 && 
b[8612] == 8612 && 
b[8613] == 8613 && 
b[8614] == 8614 && 
b[8615] == 8615 && 
b[8616] == 8616 && 
b[8617] == 8617 && 
b[8618] == 8618 && 
b[8619] == 8619 && 
b[8620] == 8620 && 
b[8621] == 8621 && 
b[8622] == 8622 && 
b[8623] == 8623 && 
b[8624] == 8624 && 
b[8625] == 8625 && 
b[8626] == 8626 && 
b[8627] == 8627 && 
b[8628] == 8628 && 
b[8629] == 8629 && 
b[8630] == 8630 && 
b[8631] == 8631 && 
b[8632] == 8632 && 
b[8633] == 8633 && 
b[8634] == 8634 && 
b[8635] == 8635 && 
b[8636] == 8636 && 
b[8637] == 8637 && 
b[8638] == 8638 && 
b[8639] == 8639 && 
b[8640] == 8640 && 
b[8641] == 8641 && 
b[8642] == 8642 && 
b[8643] == 8643 && 
b[8644] == 8644 && 
b[8645] == 8645 && 
b[8646] == 8646 && 
b[8647] == 8647 && 
b[8648] == 8648 && 
b[8649] == 8649 && 
b[8650] == 8650 && 
b[8651] == 8651 && 
b[8652] == 8652 && 
b[8653] == 8653 && 
b[8654] == 8654 && 
b[8655] == 8655 && 
b[8656] == 8656 && 
b[8657] == 8657 && 
b[8658] == 8658 && 
b[8659] == 8659 && 
b[8660] == 8660 && 
b[8661] == 8661 && 
b[8662] == 8662 && 
b[8663] == 8663 && 
b[8664] == 8664 && 
b[8665] == 8665 && 
b[8666] == 8666 && 
b[8667] == 8667 && 
b[8668] == 8668 && 
b[8669] == 8669 && 
b[8670] == 8670 && 
b[8671] == 8671 && 
b[8672] == 8672 && 
b[8673] == 8673 && 
b[8674] == 8674 && 
b[8675] == 8675 && 
b[8676] == 8676 && 
b[8677] == 8677 && 
b[8678] == 8678 && 
b[8679] == 8679 && 
b[8680] == 8680 && 
b[8681] == 8681 && 
b[8682] == 8682 && 
b[8683] == 8683 && 
b[8684] == 8684 && 
b[8685] == 8685 && 
b[8686] == 8686 && 
b[8687] == 8687 && 
b[8688] == 8688 && 
b[8689] == 8689 && 
b[8690] == 8690 && 
b[8691] == 8691 && 
b[8692] == 8692 && 
b[8693] == 8693 && 
b[8694] == 8694 && 
b[8695] == 8695 && 
b[8696] == 8696 && 
b[8697] == 8697 && 
b[8698] == 8698 && 
b[8699] == 8699 && 
b[8700] == 8700 && 
b[8701] == 8701 && 
b[8702] == 8702 && 
b[8703] == 8703 && 
b[8704] == 8704 && 
b[8705] == 8705 && 
b[8706] == 8706 && 
b[8707] == 8707 && 
b[8708] == 8708 && 
b[8709] == 8709 && 
b[8710] == 8710 && 
b[8711] == 8711 && 
b[8712] == 8712 && 
b[8713] == 8713 && 
b[8714] == 8714 && 
b[8715] == 8715 && 
b[8716] == 8716 && 
b[8717] == 8717 && 
b[8718] == 8718 && 
b[8719] == 8719 && 
b[8720] == 8720 && 
b[8721] == 8721 && 
b[8722] == 8722 && 
b[8723] == 8723 && 
b[8724] == 8724 && 
b[8725] == 8725 && 
b[8726] == 8726 && 
b[8727] == 8727 && 
b[8728] == 8728 && 
b[8729] == 8729 && 
b[8730] == 8730 && 
b[8731] == 8731 && 
b[8732] == 8732 && 
b[8733] == 8733 && 
b[8734] == 8734 && 
b[8735] == 8735 && 
b[8736] == 8736 && 
b[8737] == 8737 && 
b[8738] == 8738 && 
b[8739] == 8739 && 
b[8740] == 8740 && 
b[8741] == 8741 && 
b[8742] == 8742 && 
b[8743] == 8743 && 
b[8744] == 8744 && 
b[8745] == 8745 && 
b[8746] == 8746 && 
b[8747] == 8747 && 
b[8748] == 8748 && 
b[8749] == 8749 && 
b[8750] == 8750 && 
b[8751] == 8751 && 
b[8752] == 8752 && 
b[8753] == 8753 && 
b[8754] == 8754 && 
b[8755] == 8755 && 
b[8756] == 8756 && 
b[8757] == 8757 && 
b[8758] == 8758 && 
b[8759] == 8759 && 
b[8760] == 8760 && 
b[8761] == 8761 && 
b[8762] == 8762 && 
b[8763] == 8763 && 
b[8764] == 8764 && 
b[8765] == 8765 && 
b[8766] == 8766 && 
b[8767] == 8767 && 
b[8768] == 8768 && 
b[8769] == 8769 && 
b[8770] == 8770 && 
b[8771] == 8771 && 
b[8772] == 8772 && 
b[8773] == 8773 && 
b[8774] == 8774 && 
b[8775] == 8775 && 
b[8776] == 8776 && 
b[8777] == 8777 && 
b[8778] == 8778 && 
b[8779] == 8779 && 
b[8780] == 8780 && 
b[8781] == 8781 && 
b[8782] == 8782 && 
b[8783] == 8783 && 
b[8784] == 8784 && 
b[8785] == 8785 && 
b[8786] == 8786 && 
b[8787] == 8787 && 
b[8788] == 8788 && 
b[8789] == 8789 && 
b[8790] == 8790 && 
b[8791] == 8791 && 
b[8792] == 8792 && 
b[8793] == 8793 && 
b[8794] == 8794 && 
b[8795] == 8795 && 
b[8796] == 8796 && 
b[8797] == 8797 && 
b[8798] == 8798 && 
b[8799] == 8799 && 
b[8800] == 8800 && 
b[8801] == 8801 && 
b[8802] == 8802 && 
b[8803] == 8803 && 
b[8804] == 8804 && 
b[8805] == 8805 && 
b[8806] == 8806 && 
b[8807] == 8807 && 
b[8808] == 8808 && 
b[8809] == 8809 && 
b[8810] == 8810 && 
b[8811] == 8811 && 
b[8812] == 8812 && 
b[8813] == 8813 && 
b[8814] == 8814 && 
b[8815] == 8815 && 
b[8816] == 8816 && 
b[8817] == 8817 && 
b[8818] == 8818 && 
b[8819] == 8819 && 
b[8820] == 8820 && 
b[8821] == 8821 && 
b[8822] == 8822 && 
b[8823] == 8823 && 
b[8824] == 8824 && 
b[8825] == 8825 && 
b[8826] == 8826 && 
b[8827] == 8827 && 
b[8828] == 8828 && 
b[8829] == 8829 && 
b[8830] == 8830 && 
b[8831] == 8831 && 
b[8832] == 8832 && 
b[8833] == 8833 && 
b[8834] == 8834 && 
b[8835] == 8835 && 
b[8836] == 8836 && 
b[8837] == 8837 && 
b[8838] == 8838 && 
b[8839] == 8839 && 
b[8840] == 8840 && 
b[8841] == 8841 && 
b[8842] == 8842 && 
b[8843] == 8843 && 
b[8844] == 8844 && 
b[8845] == 8845 && 
b[8846] == 8846 && 
b[8847] == 8847 && 
b[8848] == 8848 && 
b[8849] == 8849 && 
b[8850] == 8850 && 
b[8851] == 8851 && 
b[8852] == 8852 && 
b[8853] == 8853 && 
b[8854] == 8854 && 
b[8855] == 8855 && 
b[8856] == 8856 && 
b[8857] == 8857 && 
b[8858] == 8858 && 
b[8859] == 8859 && 
b[8860] == 8860 && 
b[8861] == 8861 && 
b[8862] == 8862 && 
b[8863] == 8863 && 
b[8864] == 8864 && 
b[8865] == 8865 && 
b[8866] == 8866 && 
b[8867] == 8867 && 
b[8868] == 8868 && 
b[8869] == 8869 && 
b[8870] == 8870 && 
b[8871] == 8871 && 
b[8872] == 8872 && 
b[8873] == 8873 && 
b[8874] == 8874 && 
b[8875] == 8875 && 
b[8876] == 8876 && 
b[8877] == 8877 && 
b[8878] == 8878 && 
b[8879] == 8879 && 
b[8880] == 8880 && 
b[8881] == 8881 && 
b[8882] == 8882 && 
b[8883] == 8883 && 
b[8884] == 8884 && 
b[8885] == 8885 && 
b[8886] == 8886 && 
b[8887] == 8887 && 
b[8888] == 8888 && 
b[8889] == 8889 && 
b[8890] == 8890 && 
b[8891] == 8891 && 
b[8892] == 8892 && 
b[8893] == 8893 && 
b[8894] == 8894 && 
b[8895] == 8895 && 
b[8896] == 8896 && 
b[8897] == 8897 && 
b[8898] == 8898 && 
b[8899] == 8899 && 
b[8900] == 8900 && 
b[8901] == 8901 && 
b[8902] == 8902 && 
b[8903] == 8903 && 
b[8904] == 8904 && 
b[8905] == 8905 && 
b[8906] == 8906 && 
b[8907] == 8907 && 
b[8908] == 8908 && 
b[8909] == 8909 && 
b[8910] == 8910 && 
b[8911] == 8911 && 
b[8912] == 8912 && 
b[8913] == 8913 && 
b[8914] == 8914 && 
b[8915] == 8915 && 
b[8916] == 8916 && 
b[8917] == 8917 && 
b[8918] == 8918 && 
b[8919] == 8919 && 
b[8920] == 8920 && 
b[8921] == 8921 && 
b[8922] == 8922 && 
b[8923] == 8923 && 
b[8924] == 8924 && 
b[8925] == 8925 && 
b[8926] == 8926 && 
b[8927] == 8927 && 
b[8928] == 8928 && 
b[8929] == 8929 && 
b[8930] == 8930 && 
b[8931] == 8931 && 
b[8932] == 8932 && 
b[8933] == 8933 && 
b[8934] == 8934 && 
b[8935] == 8935 && 
b[8936] == 8936 && 
b[8937] == 8937 && 
b[8938] == 8938 && 
b[8939] == 8939 && 
b[8940] == 8940 && 
b[8941] == 8941 && 
b[8942] == 8942 && 
b[8943] == 8943 && 
b[8944] == 8944 && 
b[8945] == 8945 && 
b[8946] == 8946 && 
b[8947] == 8947 && 
b[8948] == 8948 && 
b[8949] == 8949 && 
b[8950] == 8950 && 
b[8951] == 8951 && 
b[8952] == 8952 && 
b[8953] == 8953 && 
b[8954] == 8954 && 
b[8955] == 8955 && 
b[8956] == 8956 && 
b[8957] == 8957 && 
b[8958] == 8958 && 
b[8959] == 8959 && 
b[8960] == 8960 && 
b[8961] == 8961 && 
b[8962] == 8962 && 
b[8963] == 8963 && 
b[8964] == 8964 && 
b[8965] == 8965 && 
b[8966] == 8966 && 
b[8967] == 8967 && 
b[8968] == 8968 && 
b[8969] == 8969 && 
b[8970] == 8970 && 
b[8971] == 8971 && 
b[8972] == 8972 && 
b[8973] == 8973 && 
b[8974] == 8974 && 
b[8975] == 8975 && 
b[8976] == 8976 && 
b[8977] == 8977 && 
b[8978] == 8978 && 
b[8979] == 8979 && 
b[8980] == 8980 && 
b[8981] == 8981 && 
b[8982] == 8982 && 
b[8983] == 8983 && 
b[8984] == 8984 && 
b[8985] == 8985 && 
b[8986] == 8986 && 
b[8987] == 8987 && 
b[8988] == 8988 && 
b[8989] == 8989 && 
b[8990] == 8990 && 
b[8991] == 8991 && 
b[8992] == 8992 && 
b[8993] == 8993 && 
b[8994] == 8994 && 
b[8995] == 8995 && 
b[8996] == 8996 && 
b[8997] == 8997 && 
b[8998] == 8998 && 
b[8999] == 8999 && 
b[9000] == 9000 && 
b[9001] == 9001 && 
b[9002] == 9002 && 
b[9003] == 9003 && 
b[9004] == 9004 && 
b[9005] == 9005 && 
b[9006] == 9006 && 
b[9007] == 9007 && 
b[9008] == 9008 && 
b[9009] == 9009 && 
b[9010] == 9010 && 
b[9011] == 9011 && 
b[9012] == 9012 && 
b[9013] == 9013 && 
b[9014] == 9014 && 
b[9015] == 9015 && 
b[9016] == 9016 && 
b[9017] == 9017 && 
b[9018] == 9018 && 
b[9019] == 9019 && 
b[9020] == 9020 && 
b[9021] == 9021 && 
b[9022] == 9022 && 
b[9023] == 9023 && 
b[9024] == 9024 && 
b[9025] == 9025 && 
b[9026] == 9026 && 
b[9027] == 9027 && 
b[9028] == 9028 && 
b[9029] == 9029 && 
b[9030] == 9030 && 
b[9031] == 9031 && 
b[9032] == 9032 && 
b[9033] == 9033 && 
b[9034] == 9034 && 
b[9035] == 9035 && 
b[9036] == 9036 && 
b[9037] == 9037 && 
b[9038] == 9038 && 
b[9039] == 9039 && 
b[9040] == 9040 && 
b[9041] == 9041 && 
b[9042] == 9042 && 
b[9043] == 9043 && 
b[9044] == 9044 && 
b[9045] == 9045 && 
b[9046] == 9046 && 
b[9047] == 9047 && 
b[9048] == 9048 && 
b[9049] == 9049 && 
b[9050] == 9050 && 
b[9051] == 9051 && 
b[9052] == 9052 && 
b[9053] == 9053 && 
b[9054] == 9054 && 
b[9055] == 9055 && 
b[9056] == 9056 && 
b[9057] == 9057 && 
b[9058] == 9058 && 
b[9059] == 9059 && 
b[9060] == 9060 && 
b[9061] == 9061 && 
b[9062] == 9062 && 
b[9063] == 9063 && 
b[9064] == 9064 && 
b[9065] == 9065 && 
b[9066] == 9066 && 
b[9067] == 9067 && 
b[9068] == 9068 && 
b[9069] == 9069 && 
b[9070] == 9070 && 
b[9071] == 9071 && 
b[9072] == 9072 && 
b[9073] == 9073 && 
b[9074] == 9074 && 
b[9075] == 9075 && 
b[9076] == 9076 && 
b[9077] == 9077 && 
b[9078] == 9078 && 
b[9079] == 9079 && 
b[9080] == 9080 && 
b[9081] == 9081 && 
b[9082] == 9082 && 
b[9083] == 9083 && 
b[9084] == 9084 && 
b[9085] == 9085 && 
b[9086] == 9086 && 
b[9087] == 9087 && 
b[9088] == 9088 && 
b[9089] == 9089 && 
b[9090] == 9090 && 
b[9091] == 9091 && 
b[9092] == 9092 && 
b[9093] == 9093 && 
b[9094] == 9094 && 
b[9095] == 9095 && 
b[9096] == 9096 && 
b[9097] == 9097 && 
b[9098] == 9098 && 
b[9099] == 9099 && 
b[9100] == 9100 && 
b[9101] == 9101 && 
b[9102] == 9102 && 
b[9103] == 9103 && 
b[9104] == 9104 && 
b[9105] == 9105 && 
b[9106] == 9106 && 
b[9107] == 9107 && 
b[9108] == 9108 && 
b[9109] == 9109 && 
b[9110] == 9110 && 
b[9111] == 9111 && 
b[9112] == 9112 && 
b[9113] == 9113 && 
b[9114] == 9114 && 
b[9115] == 9115 && 
b[9116] == 9116 && 
b[9117] == 9117 && 
b[9118] == 9118 && 
b[9119] == 9119 && 
b[9120] == 9120 && 
b[9121] == 9121 && 
b[9122] == 9122 && 
b[9123] == 9123 && 
b[9124] == 9124 && 
b[9125] == 9125 && 
b[9126] == 9126 && 
b[9127] == 9127 && 
b[9128] == 9128 && 
b[9129] == 9129 && 
b[9130] == 9130 && 
b[9131] == 9131 && 
b[9132] == 9132 && 
b[9133] == 9133 && 
b[9134] == 9134 && 
b[9135] == 9135 && 
b[9136] == 9136 && 
b[9137] == 9137 && 
b[9138] == 9138 && 
b[9139] == 9139 && 
b[9140] == 9140 && 
b[9141] == 9141 && 
b[9142] == 9142 && 
b[9143] == 9143 && 
b[9144] == 9144 && 
b[9145] == 9145 && 
b[9146] == 9146 && 
b[9147] == 9147 && 
b[9148] == 9148 && 
b[9149] == 9149 && 
b[9150] == 9150 && 
b[9151] == 9151 && 
b[9152] == 9152 && 
b[9153] == 9153 && 
b[9154] == 9154 && 
b[9155] == 9155 && 
b[9156] == 9156 && 
b[9157] == 9157 && 
b[9158] == 9158 && 
b[9159] == 9159 && 
b[9160] == 9160 && 
b[9161] == 9161 && 
b[9162] == 9162 && 
b[9163] == 9163 && 
b[9164] == 9164 && 
b[9165] == 9165 && 
b[9166] == 9166 && 
b[9167] == 9167 && 
b[9168] == 9168 && 
b[9169] == 9169 && 
b[9170] == 9170 && 
b[9171] == 9171 && 
b[9172] == 9172 && 
b[9173] == 9173 && 
b[9174] == 9174 && 
b[9175] == 9175 && 
b[9176] == 9176 && 
b[9177] == 9177 && 
b[9178] == 9178 && 
b[9179] == 9179 && 
b[9180] == 9180 && 
b[9181] == 9181 && 
b[9182] == 9182 && 
b[9183] == 9183 && 
b[9184] == 9184 && 
b[9185] == 9185 && 
b[9186] == 9186 && 
b[9187] == 9187 && 
b[9188] == 9188 && 
b[9189] == 9189 && 
b[9190] == 9190 && 
b[9191] == 9191 && 
b[9192] == 9192 && 
b[9193] == 9193 && 
b[9194] == 9194 && 
b[9195] == 9195 && 
b[9196] == 9196 && 
b[9197] == 9197 && 
b[9198] == 9198 && 
b[9199] == 9199 && 
b[9200] == 9200 && 
b[9201] == 9201 && 
b[9202] == 9202 && 
b[9203] == 9203 && 
b[9204] == 9204 && 
b[9205] == 9205 && 
b[9206] == 9206 && 
b[9207] == 9207 && 
b[9208] == 9208 && 
b[9209] == 9209 && 
b[9210] == 9210 && 
b[9211] == 9211 && 
b[9212] == 9212 && 
b[9213] == 9213 && 
b[9214] == 9214 && 
b[9215] == 9215 && 
b[9216] == 9216 && 
b[9217] == 9217 && 
b[9218] == 9218 && 
b[9219] == 9219 && 
b[9220] == 9220 && 
b[9221] == 9221 && 
b[9222] == 9222 && 
b[9223] == 9223 && 
b[9224] == 9224 && 
b[9225] == 9225 && 
b[9226] == 9226 && 
b[9227] == 9227 && 
b[9228] == 9228 && 
b[9229] == 9229 && 
b[9230] == 9230 && 
b[9231] == 9231 && 
b[9232] == 9232 && 
b[9233] == 9233 && 
b[9234] == 9234 && 
b[9235] == 9235 && 
b[9236] == 9236 && 
b[9237] == 9237 && 
b[9238] == 9238 && 
b[9239] == 9239 && 
b[9240] == 9240 && 
b[9241] == 9241 && 
b[9242] == 9242 && 
b[9243] == 9243 && 
b[9244] == 9244 && 
b[9245] == 9245 && 
b[9246] == 9246 && 
b[9247] == 9247 && 
b[9248] == 9248 && 
b[9249] == 9249 && 
b[9250] == 9250 && 
b[9251] == 9251 && 
b[9252] == 9252 && 
b[9253] == 9253 && 
b[9254] == 9254 && 
b[9255] == 9255 && 
b[9256] == 9256 && 
b[9257] == 9257 && 
b[9258] == 9258 && 
b[9259] == 9259 && 
b[9260] == 9260 && 
b[9261] == 9261 && 
b[9262] == 9262 && 
b[9263] == 9263 && 
b[9264] == 9264 && 
b[9265] == 9265 && 
b[9266] == 9266 && 
b[9267] == 9267 && 
b[9268] == 9268 && 
b[9269] == 9269 && 
b[9270] == 9270 && 
b[9271] == 9271 && 
b[9272] == 9272 && 
b[9273] == 9273 && 
b[9274] == 9274 && 
b[9275] == 9275 && 
b[9276] == 9276 && 
b[9277] == 9277 && 
b[9278] == 9278 && 
b[9279] == 9279 && 
b[9280] == 9280 && 
b[9281] == 9281 && 
b[9282] == 9282 && 
b[9283] == 9283 && 
b[9284] == 9284 && 
b[9285] == 9285 && 
b[9286] == 9286 && 
b[9287] == 9287 && 
b[9288] == 9288 && 
b[9289] == 9289 && 
b[9290] == 9290 && 
b[9291] == 9291 && 
b[9292] == 9292 && 
b[9293] == 9293 && 
b[9294] == 9294 && 
b[9295] == 9295 && 
b[9296] == 9296 && 
b[9297] == 9297 && 
b[9298] == 9298 && 
b[9299] == 9299 && 
b[9300] == 9300 && 
b[9301] == 9301 && 
b[9302] == 9302 && 
b[9303] == 9303 && 
b[9304] == 9304 && 
b[9305] == 9305 && 
b[9306] == 9306 && 
b[9307] == 9307 && 
b[9308] == 9308 && 
b[9309] == 9309 && 
b[9310] == 9310 && 
b[9311] == 9311 && 
b[9312] == 9312 && 
b[9313] == 9313 && 
b[9314] == 9314 && 
b[9315] == 9315 && 
b[9316] == 9316 && 
b[9317] == 9317 && 
b[9318] == 9318 && 
b[9319] == 9319 && 
b[9320] == 9320 && 
b[9321] == 9321 && 
b[9322] == 9322 && 
b[9323] == 9323 && 
b[9324] == 9324 && 
b[9325] == 9325 && 
b[9326] == 9326 && 
b[9327] == 9327 && 
b[9328] == 9328 && 
b[9329] == 9329 && 
b[9330] == 9330 && 
b[9331] == 9331 && 
b[9332] == 9332 && 
b[9333] == 9333 && 
b[9334] == 9334 && 
b[9335] == 9335 && 
b[9336] == 9336 && 
b[9337] == 9337 && 
b[9338] == 9338 && 
b[9339] == 9339 && 
b[9340] == 9340 && 
b[9341] == 9341 && 
b[9342] == 9342 && 
b[9343] == 9343 && 
b[9344] == 9344 && 
b[9345] == 9345 && 
b[9346] == 9346 && 
b[9347] == 9347 && 
b[9348] == 9348 && 
b[9349] == 9349 && 
b[9350] == 9350 && 
b[9351] == 9351 && 
b[9352] == 9352 && 
b[9353] == 9353 && 
b[9354] == 9354 && 
b[9355] == 9355 && 
b[9356] == 9356 && 
b[9357] == 9357 && 
b[9358] == 9358 && 
b[9359] == 9359 && 
b[9360] == 9360 && 
b[9361] == 9361 && 
b[9362] == 9362 && 
b[9363] == 9363 && 
b[9364] == 9364 && 
b[9365] == 9365 && 
b[9366] == 9366 && 
b[9367] == 9367 && 
b[9368] == 9368 && 
b[9369] == 9369 && 
b[9370] == 9370 && 
b[9371] == 9371 && 
b[9372] == 9372 && 
b[9373] == 9373 && 
b[9374] == 9374 && 
b[9375] == 9375 && 
b[9376] == 9376 && 
b[9377] == 9377 && 
b[9378] == 9378 && 
b[9379] == 9379 && 
b[9380] == 9380 && 
b[9381] == 9381 && 
b[9382] == 9382 && 
b[9383] == 9383 && 
b[9384] == 9384 && 
b[9385] == 9385 && 
b[9386] == 9386 && 
b[9387] == 9387 && 
b[9388] == 9388 && 
b[9389] == 9389 && 
b[9390] == 9390 && 
b[9391] == 9391 && 
b[9392] == 9392 && 
b[9393] == 9393 && 
b[9394] == 9394 && 
b[9395] == 9395 && 
b[9396] == 9396 && 
b[9397] == 9397 && 
b[9398] == 9398 && 
b[9399] == 9399 && 
b[9400] == 9400 && 
b[9401] == 9401 && 
b[9402] == 9402 && 
b[9403] == 9403 && 
b[9404] == 9404 && 
b[9405] == 9405 && 
b[9406] == 9406 && 
b[9407] == 9407 && 
b[9408] == 9408 && 
b[9409] == 9409 && 
b[9410] == 9410 && 
b[9411] == 9411 && 
b[9412] == 9412 && 
b[9413] == 9413 && 
b[9414] == 9414 && 
b[9415] == 9415 && 
b[9416] == 9416 && 
b[9417] == 9417 && 
b[9418] == 9418 && 
b[9419] == 9419 && 
b[9420] == 9420 && 
b[9421] == 9421 && 
b[9422] == 9422 && 
b[9423] == 9423 && 
b[9424] == 9424 && 
b[9425] == 9425 && 
b[9426] == 9426 && 
b[9427] == 9427 && 
b[9428] == 9428 && 
b[9429] == 9429 && 
b[9430] == 9430 && 
b[9431] == 9431 && 
b[9432] == 9432 && 
b[9433] == 9433 && 
b[9434] == 9434 && 
b[9435] == 9435 && 
b[9436] == 9436 && 
b[9437] == 9437 && 
b[9438] == 9438 && 
b[9439] == 9439 && 
b[9440] == 9440 && 
b[9441] == 9441 && 
b[9442] == 9442 && 
b[9443] == 9443 && 
b[9444] == 9444 && 
b[9445] == 9445 && 
b[9446] == 9446 && 
b[9447] == 9447 && 
b[9448] == 9448 && 
b[9449] == 9449 && 
b[9450] == 9450 && 
b[9451] == 9451 && 
b[9452] == 9452 && 
b[9453] == 9453 && 
b[9454] == 9454 && 
b[9455] == 9455 && 
b[9456] == 9456 && 
b[9457] == 9457 && 
b[9458] == 9458 && 
b[9459] == 9459 && 
b[9460] == 9460 && 
b[9461] == 9461 && 
b[9462] == 9462 && 
b[9463] == 9463 && 
b[9464] == 9464 && 
b[9465] == 9465 && 
b[9466] == 9466 && 
b[9467] == 9467 && 
b[9468] == 9468 && 
b[9469] == 9469 && 
b[9470] == 9470 && 
b[9471] == 9471 && 
b[9472] == 9472 && 
b[9473] == 9473 && 
b[9474] == 9474 && 
b[9475] == 9475 && 
b[9476] == 9476 && 
b[9477] == 9477 && 
b[9478] == 9478 && 
b[9479] == 9479 && 
b[9480] == 9480 && 
b[9481] == 9481 && 
b[9482] == 9482 && 
b[9483] == 9483 && 
b[9484] == 9484 && 
b[9485] == 9485 && 
b[9486] == 9486 && 
b[9487] == 9487 && 
b[9488] == 9488 && 
b[9489] == 9489 && 
b[9490] == 9490 && 
b[9491] == 9491 && 
b[9492] == 9492 && 
b[9493] == 9493 && 
b[9494] == 9494 && 
b[9495] == 9495 && 
b[9496] == 9496 && 
b[9497] == 9497 && 
b[9498] == 9498 && 
b[9499] == 9499 && 
b[9500] == 9500 && 
b[9501] == 9501 && 
b[9502] == 9502 && 
b[9503] == 9503 && 
b[9504] == 9504 && 
b[9505] == 9505 && 
b[9506] == 9506 && 
b[9507] == 9507 && 
b[9508] == 9508 && 
b[9509] == 9509 && 
b[9510] == 9510 && 
b[9511] == 9511 && 
b[9512] == 9512 && 
b[9513] == 9513 && 
b[9514] == 9514 && 
b[9515] == 9515 && 
b[9516] == 9516 && 
b[9517] == 9517 && 
b[9518] == 9518 && 
b[9519] == 9519 && 
b[9520] == 9520 && 
b[9521] == 9521 && 
b[9522] == 9522 && 
b[9523] == 9523 && 
b[9524] == 9524 && 
b[9525] == 9525 && 
b[9526] == 9526 && 
b[9527] == 9527 && 
b[9528] == 9528 && 
b[9529] == 9529 && 
b[9530] == 9530 && 
b[9531] == 9531 && 
b[9532] == 9532 && 
b[9533] == 9533 && 
b[9534] == 9534 && 
b[9535] == 9535 && 
b[9536] == 9536 && 
b[9537] == 9537 && 
b[9538] == 9538 && 
b[9539] == 9539 && 
b[9540] == 9540 && 
b[9541] == 9541 && 
b[9542] == 9542 && 
b[9543] == 9543 && 
b[9544] == 9544 && 
b[9545] == 9545 && 
b[9546] == 9546 && 
b[9547] == 9547 && 
b[9548] == 9548 && 
b[9549] == 9549 && 
b[9550] == 9550 && 
b[9551] == 9551 && 
b[9552] == 9552 && 
b[9553] == 9553 && 
b[9554] == 9554 && 
b[9555] == 9555 && 
b[9556] == 9556 && 
b[9557] == 9557 && 
b[9558] == 9558 && 
b[9559] == 9559 && 
b[9560] == 9560 && 
b[9561] == 9561 && 
b[9562] == 9562 && 
b[9563] == 9563 && 
b[9564] == 9564 && 
b[9565] == 9565 && 
b[9566] == 9566 && 
b[9567] == 9567 && 
b[9568] == 9568 && 
b[9569] == 9569 && 
b[9570] == 9570 && 
b[9571] == 9571 && 
b[9572] == 9572 && 
b[9573] == 9573 && 
b[9574] == 9574 && 
b[9575] == 9575 && 
b[9576] == 9576 && 
b[9577] == 9577 && 
b[9578] == 9578 && 
b[9579] == 9579 && 
b[9580] == 9580 && 
b[9581] == 9581 && 
b[9582] == 9582 && 
b[9583] == 9583 && 
b[9584] == 9584 && 
b[9585] == 9585 && 
b[9586] == 9586 && 
b[9587] == 9587 && 
b[9588] == 9588 && 
b[9589] == 9589 && 
b[9590] == 9590 && 
b[9591] == 9591 && 
b[9592] == 9592 && 
b[9593] == 9593 && 
b[9594] == 9594 && 
b[9595] == 9595 && 
b[9596] == 9596 && 
b[9597] == 9597 && 
b[9598] == 9598 && 
b[9599] == 9599 && 
b[9600] == 9600 && 
b[9601] == 9601 && 
b[9602] == 9602 && 
b[9603] == 9603 && 
b[9604] == 9604 && 
b[9605] == 9605 && 
b[9606] == 9606 && 
b[9607] == 9607 && 
b[9608] == 9608 && 
b[9609] == 9609 && 
b[9610] == 9610 && 
b[9611] == 9611 && 
b[9612] == 9612 && 
b[9613] == 9613 && 
b[9614] == 9614 && 
b[9615] == 9615 && 
b[9616] == 9616 && 
b[9617] == 9617 && 
b[9618] == 9618 && 
b[9619] == 9619 && 
b[9620] == 9620 && 
b[9621] == 9621 && 
b[9622] == 9622 && 
b[9623] == 9623 && 
b[9624] == 9624 && 
b[9625] == 9625 && 
b[9626] == 9626 && 
b[9627] == 9627 && 
b[9628] == 9628 && 
b[9629] == 9629 && 
b[9630] == 9630 && 
b[9631] == 9631 && 
b[9632] == 9632 && 
b[9633] == 9633 && 
b[9634] == 9634 && 
b[9635] == 9635 && 
b[9636] == 9636 && 
b[9637] == 9637 && 
b[9638] == 9638 && 
b[9639] == 9639 && 
b[9640] == 9640 && 
b[9641] == 9641 && 
b[9642] == 9642 && 
b[9643] == 9643 && 
b[9644] == 9644 && 
b[9645] == 9645 && 
b[9646] == 9646 && 
b[9647] == 9647 && 
b[9648] == 9648 && 
b[9649] == 9649 && 
b[9650] == 9650 && 
b[9651] == 9651 && 
b[9652] == 9652 && 
b[9653] == 9653 && 
b[9654] == 9654 && 
b[9655] == 9655 && 
b[9656] == 9656 && 
b[9657] == 9657 && 
b[9658] == 9658 && 
b[9659] == 9659 && 
b[9660] == 9660 && 
b[9661] == 9661 && 
b[9662] == 9662 && 
b[9663] == 9663 && 
b[9664] == 9664 && 
b[9665] == 9665 && 
b[9666] == 9666 && 
b[9667] == 9667 && 
b[9668] == 9668 && 
b[9669] == 9669 && 
b[9670] == 9670 && 
b[9671] == 9671 && 
b[9672] == 9672 && 
b[9673] == 9673 && 
b[9674] == 9674 && 
b[9675] == 9675 && 
b[9676] == 9676 && 
b[9677] == 9677 && 
b[9678] == 9678 && 
b[9679] == 9679 && 
b[9680] == 9680 && 
b[9681] == 9681 && 
b[9682] == 9682 && 
b[9683] == 9683 && 
b[9684] == 9684 && 
b[9685] == 9685 && 
b[9686] == 9686 && 
b[9687] == 9687 && 
b[9688] == 9688 && 
b[9689] == 9689 && 
b[9690] == 9690 && 
b[9691] == 9691 && 
b[9692] == 9692 && 
b[9693] == 9693 && 
b[9694] == 9694 && 
b[9695] == 9695 && 
b[9696] == 9696 && 
b[9697] == 9697 && 
b[9698] == 9698 && 
b[9699] == 9699 && 
b[9700] == 9700 && 
b[9701] == 9701 && 
b[9702] == 9702 && 
b[9703] == 9703 && 
b[9704] == 9704 && 
b[9705] == 9705 && 
b[9706] == 9706 && 
b[9707] == 9707 && 
b[9708] == 9708 && 
b[9709] == 9709 && 
b[9710] == 9710 && 
b[9711] == 9711 && 
b[9712] == 9712 && 
b[9713] == 9713 && 
b[9714] == 9714 && 
b[9715] == 9715 && 
b[9716] == 9716 && 
b[9717] == 9717 && 
b[9718] == 9718 && 
b[9719] == 9719 && 
b[9720] == 9720 && 
b[9721] == 9721 && 
b[9722] == 9722 && 
b[9723] == 9723 && 
b[9724] == 9724 && 
b[9725] == 9725 && 
b[9726] == 9726 && 
b[9727] == 9727 && 
b[9728] == 9728 && 
b[9729] == 9729 && 
b[9730] == 9730 && 
b[9731] == 9731 && 
b[9732] == 9732 && 
b[9733] == 9733 && 
b[9734] == 9734 && 
b[9735] == 9735 && 
b[9736] == 9736 && 
b[9737] == 9737 && 
b[9738] == 9738 && 
b[9739] == 9739 && 
b[9740] == 9740 && 
b[9741] == 9741 && 
b[9742] == 9742 && 
b[9743] == 9743 && 
b[9744] == 9744 && 
b[9745] == 9745 && 
b[9746] == 9746 && 
b[9747] == 9747 && 
b[9748] == 9748 && 
b[9749] == 9749 && 
b[9750] == 9750 && 
b[9751] == 9751 && 
b[9752] == 9752 && 
b[9753] == 9753 && 
b[9754] == 9754 && 
b[9755] == 9755 && 
b[9756] == 9756 && 
b[9757] == 9757 && 
b[9758] == 9758 && 
b[9759] == 9759 && 
b[9760] == 9760 && 
b[9761] == 9761 && 
b[9762] == 9762 && 
b[9763] == 9763 && 
b[9764] == 9764 && 
b[9765] == 9765 && 
b[9766] == 9766 && 
b[9767] == 9767 && 
b[9768] == 9768 && 
b[9769] == 9769 && 
b[9770] == 9770 && 
b[9771] == 9771 && 
b[9772] == 9772 && 
b[9773] == 9773 && 
b[9774] == 9774 && 
b[9775] == 9775 && 
b[9776] == 9776 && 
b[9777] == 9777 && 
b[9778] == 9778 && 
b[9779] == 9779 && 
b[9780] == 9780 && 
b[9781] == 9781 && 
b[9782] == 9782 && 
b[9783] == 9783 && 
b[9784] == 9784 && 
b[9785] == 9785 && 
b[9786] == 9786 && 
b[9787] == 9787 && 
b[9788] == 9788 && 
b[9789] == 9789 && 
b[9790] == 9790 && 
b[9791] == 9791 && 
b[9792] == 9792 && 
b[9793] == 9793 && 
b[9794] == 9794 && 
b[9795] == 9795 && 
b[9796] == 9796 && 
b[9797] == 9797 && 
b[9798] == 9798 && 
b[9799] == 9799 && 
b[9800] == 9800 && 
b[9801] == 9801 && 
b[9802] == 9802 && 
b[9803] == 9803 && 
b[9804] == 9804 && 
b[9805] == 9805 && 
b[9806] == 9806 && 
b[9807] == 9807 && 
b[9808] == 9808 && 
b[9809] == 9809 && 
b[9810] == 9810 && 
b[9811] == 9811 && 
b[9812] == 9812 && 
b[9813] == 9813 && 
b[9814] == 9814 && 
b[9815] == 9815 && 
b[9816] == 9816 && 
b[9817] == 9817 && 
b[9818] == 9818 && 
b[9819] == 9819 && 
b[9820] == 9820 && 
b[9821] == 9821 && 
b[9822] == 9822 && 
b[9823] == 9823 && 
b[9824] == 9824 && 
b[9825] == 9825 && 
b[9826] == 9826 && 
b[9827] == 9827 && 
b[9828] == 9828 && 
b[9829] == 9829 && 
b[9830] == 9830 && 
b[9831] == 9831 && 
b[9832] == 9832 && 
b[9833] == 9833 && 
b[9834] == 9834 && 
b[9835] == 9835 && 
b[9836] == 9836 && 
b[9837] == 9837 && 
b[9838] == 9838 && 
b[9839] == 9839 && 
b[9840] == 9840 && 
b[9841] == 9841 && 
b[9842] == 9842 && 
b[9843] == 9843 && 
b[9844] == 9844 && 
b[9845] == 9845 && 
b[9846] == 9846 && 
b[9847] == 9847 && 
b[9848] == 9848 && 
b[9849] == 9849 && 
b[9850] == 9850 && 
b[9851] == 9851 && 
b[9852] == 9852 && 
b[9853] == 9853 && 
b[9854] == 9854 && 
b[9855] == 9855 && 
b[9856] == 9856 && 
b[9857] == 9857 && 
b[9858] == 9858 && 
b[9859] == 9859 && 
b[9860] == 9860 && 
b[9861] == 9861 && 
b[9862] == 9862 && 
b[9863] == 9863 && 
b[9864] == 9864 && 
b[9865] == 9865 && 
b[9866] == 9866 && 
b[9867] == 9867 && 
b[9868] == 9868 && 
b[9869] == 9869 && 
b[9870] == 9870 && 
b[9871] == 9871 && 
b[9872] == 9872 && 
b[9873] == 9873 && 
b[9874] == 9874 && 
b[9875] == 9875 && 
b[9876] == 9876 && 
b[9877] == 9877 && 
b[9878] == 9878 && 
b[9879] == 9879 && 
b[9880] == 9880 && 
b[9881] == 9881 && 
b[9882] == 9882 && 
b[9883] == 9883 && 
b[9884] == 9884 && 
b[9885] == 9885 && 
b[9886] == 9886 && 
b[9887] == 9887 && 
b[9888] == 9888 && 
b[9889] == 9889 && 
b[9890] == 9890 && 
b[9891] == 9891 && 
b[9892] == 9892 && 
b[9893] == 9893 && 
b[9894] == 9894 && 
b[9895] == 9895 && 
b[9896] == 9896 && 
b[9897] == 9897 && 
b[9898] == 9898 && 
b[9899] == 9899 && 
b[9900] == 9900 && 
b[9901] == 9901 && 
b[9902] == 9902 && 
b[9903] == 9903 && 
b[9904] == 9904 && 
b[9905] == 9905 && 
b[9906] == 9906 && 
b[9907] == 9907 && 
b[9908] == 9908 && 
b[9909] == 9909 && 
b[9910] == 9910 && 
b[9911] == 9911 && 
b[9912] == 9912 && 
b[9913] == 9913 && 
b[9914] == 9914 && 
b[9915] == 9915 && 
b[9916] == 9916 && 
b[9917] == 9917 && 
b[9918] == 9918 && 
b[9919] == 9919 && 
b[9920] == 9920 && 
b[9921] == 9921 && 
b[9922] == 9922 && 
b[9923] == 9923 && 
b[9924] == 9924 && 
b[9925] == 9925 && 
b[9926] == 9926 && 
b[9927] == 9927 && 
b[9928] == 9928 && 
b[9929] == 9929 && 
b[9930] == 9930 && 
b[9931] == 9931 && 
b[9932] == 9932 && 
b[9933] == 9933 && 
b[9934] == 9934 && 
b[9935] == 9935 && 
b[9936] == 9936 && 
b[9937] == 9937 && 
b[9938] == 9938 && 
b[9939] == 9939 && 
b[9940] == 9940 && 
b[9941] == 9941 && 
b[9942] == 9942 && 
b[9943] == 9943 && 
b[9944] == 9944 && 
b[9945] == 9945 && 
b[9946] == 9946 && 
b[9947] == 9947 && 
b[9948] == 9948 && 
b[9949] == 9949 && 
b[9950] == 9950 && 
b[9951] == 9951 && 
b[9952] == 9952 && 
b[9953] == 9953 && 
b[9954] == 9954 && 
b[9955] == 9955 && 
b[9956] == 9956 && 
b[9957] == 9957 && 
b[9958] == 9958 && 
b[9959] == 9959 && 
b[9960] == 9960 && 
b[9961] == 9961 && 
b[9962] == 9962 && 
b[9963] == 9963 && 
b[9964] == 9964 && 
b[9965] == 9965 && 
b[9966] == 9966 && 
b[9967] == 9967 && 
b[9968] == 9968 && 
b[9969] == 9969 && 
b[9970] == 9970 && 
b[9971] == 9971 && 
b[9972] == 9972 && 
b[9973] == 9973 && 
b[9974] == 9974 && 
b[9975] == 9975 && 
b[9976] == 9976 && 
b[9977] == 9977 && 
b[9978] == 9978 && 
b[9979] == 9979 && 
b[9980] == 9980 && 
b[9981] == 9981 && 
b[9982] == 9982 && 
b[9983] == 9983 && 
b[9984] == 9984 && 
b[9985] == 9985 && 
b[9986] == 9986 && 
b[9987] == 9987 && 
b[9988] == 9988 && 
b[9989] == 9989 && 
b[9990] == 9990 && 
b[9991] == 9991 && 
b[9992] == 9992 && 
b[9993] == 9993 && 
b[9994] == 9994 && 
b[9995] == 9995 && 
b[9996] == 9996 && 
b[9997] == 9997 && 
b[9998] == 9998 && 
b[9999] == 9999 && 
b[10000] == 10000 && 
b[10001] == 10001 && 
b[10002] == 10002 && 
b[10003] == 10003 && 
b[10004] == 10004 && 
b[10005] == 10005 && 
b[10006] == 10006 && 
b[10007] == 10007 && 
b[10008] == 10008 && 
b[10009] == 10009 && 
b[10010] == 10010 && 
b[10011] == 10011 && 
b[10012] == 10012 && 
b[10013] == 10013 && 
b[10014] == 10014 && 
b[10015] == 10015 && 
b[10016] == 10016 && 
b[10017] == 10017 && 
b[10018] == 10018 && 
b[10019] == 10019 && 
b[10020] == 10020 && 
b[10021] == 10021 && 
b[10022] == 10022 && 
b[10023] == 10023 && 
b[10024] == 10024 && 
b[10025] == 10025 && 
b[10026] == 10026 && 
b[10027] == 10027 && 
b[10028] == 10028 && 
b[10029] == 10029 && 
b[10030] == 10030 && 
b[10031] == 10031 && 
b[10032] == 10032 && 
b[10033] == 10033 && 
b[10034] == 10034 && 
b[10035] == 10035 && 
b[10036] == 10036 && 
b[10037] == 10037 && 
b[10038] == 10038 && 
b[10039] == 10039 && 
b[10040] == 10040 && 
b[10041] == 10041 && 
b[10042] == 10042 && 
b[10043] == 10043 && 
b[10044] == 10044 && 
b[10045] == 10045 && 
b[10046] == 10046 && 
b[10047] == 10047 && 
b[10048] == 10048 && 
b[10049] == 10049 && 
b[10050] == 10050 && 
b[10051] == 10051 && 
b[10052] == 10052 && 
b[10053] == 10053 && 
b[10054] == 10054 && 
b[10055] == 10055 && 
b[10056] == 10056 && 
b[10057] == 10057 && 
b[10058] == 10058 && 
b[10059] == 10059 && 
b[10060] == 10060 && 
b[10061] == 10061 && 
b[10062] == 10062 && 
b[10063] == 10063 && 
b[10064] == 10064 && 
b[10065] == 10065 && 
b[10066] == 10066 && 
b[10067] == 10067 && 
b[10068] == 10068 && 
b[10069] == 10069 && 
b[10070] == 10070 && 
b[10071] == 10071 && 
b[10072] == 10072 && 
b[10073] == 10073 && 
b[10074] == 10074 && 
b[10075] == 10075 && 
b[10076] == 10076 && 
b[10077] == 10077 && 
b[10078] == 10078 && 
b[10079] == 10079 && 
b[10080] == 10080 && 
b[10081] == 10081 && 
b[10082] == 10082 && 
b[10083] == 10083 && 
b[10084] == 10084 && 
b[10085] == 10085 && 
b[10086] == 10086 && 
b[10087] == 10087 && 
b[10088] == 10088 && 
b[10089] == 10089 && 
b[10090] == 10090 && 
b[10091] == 10091 && 
b[10092] == 10092 && 
b[10093] == 10093 && 
b[10094] == 10094 && 
b[10095] == 10095 && 
b[10096] == 10096 && 
b[10097] == 10097 && 
b[10098] == 10098 && 
b[10099] == 10099 && 
b[10100] == 10100 && 
b[10101] == 10101 && 
b[10102] == 10102 && 
b[10103] == 10103 && 
b[10104] == 10104 && 
b[10105] == 10105 && 
b[10106] == 10106 && 
b[10107] == 10107 && 
b[10108] == 10108 && 
b[10109] == 10109 && 
b[10110] == 10110 && 
b[10111] == 10111 && 
b[10112] == 10112 && 
b[10113] == 10113 && 
b[10114] == 10114 && 
b[10115] == 10115 && 
b[10116] == 10116 && 
b[10117] == 10117 && 
b[10118] == 10118 && 
b[10119] == 10119 && 
b[10120] == 10120 && 
b[10121] == 10121 && 
b[10122] == 10122 && 
b[10123] == 10123 && 
b[10124] == 10124 && 
b[10125] == 10125 && 
b[10126] == 10126 && 
b[10127] == 10127 && 
b[10128] == 10128 && 
b[10129] == 10129 && 
b[10130] == 10130 && 
b[10131] == 10131 && 
b[10132] == 10132 && 
b[10133] == 10133 && 
b[10134] == 10134 && 
b[10135] == 10135 && 
b[10136] == 10136 && 
b[10137] == 10137 && 
b[10138] == 10138 && 
b[10139] == 10139 && 
b[10140] == 10140 && 
b[10141] == 10141 && 
b[10142] == 10142 && 
b[10143] == 10143 && 
b[10144] == 10144 && 
b[10145] == 10145 && 
b[10146] == 10146 && 
b[10147] == 10147 && 
b[10148] == 10148 && 
b[10149] == 10149 && 
b[10150] == 10150 && 
b[10151] == 10151 && 
b[10152] == 10152 && 
b[10153] == 10153 && 
b[10154] == 10154 && 
b[10155] == 10155 && 
b[10156] == 10156 && 
b[10157] == 10157 && 
b[10158] == 10158 && 
b[10159] == 10159 && 
b[10160] == 10160 && 
b[10161] == 10161 && 
b[10162] == 10162 && 
b[10163] == 10163 && 
b[10164] == 10164 && 
b[10165] == 10165 && 
b[10166] == 10166 && 
b[10167] == 10167 && 
b[10168] == 10168 && 
b[10169] == 10169 && 
b[10170] == 10170 && 
b[10171] == 10171 && 
b[10172] == 10172 && 
b[10173] == 10173 && 
b[10174] == 10174 && 
b[10175] == 10175 && 
b[10176] == 10176 && 
b[10177] == 10177 && 
b[10178] == 10178 && 
b[10179] == 10179 && 
b[10180] == 10180 && 
b[10181] == 10181 && 
b[10182] == 10182 && 
b[10183] == 10183 && 
b[10184] == 10184 && 
b[10185] == 10185 && 
b[10186] == 10186 && 
b[10187] == 10187 && 
b[10188] == 10188 && 
b[10189] == 10189 && 
b[10190] == 10190 && 
b[10191] == 10191 && 
b[10192] == 10192 && 
b[10193] == 10193 && 
b[10194] == 10194 && 
b[10195] == 10195 && 
b[10196] == 10196 && 
b[10197] == 10197 && 
b[10198] == 10198 && 
b[10199] == 10199 && 
b[10200] == 10200 && 
b[10201] == 10201 && 
b[10202] == 10202 && 
b[10203] == 10203 && 
b[10204] == 10204 && 
b[10205] == 10205 && 
b[10206] == 10206 && 
b[10207] == 10207 && 
b[10208] == 10208 && 
b[10209] == 10209 && 
b[10210] == 10210 && 
b[10211] == 10211 && 
b[10212] == 10212 && 
b[10213] == 10213 && 
b[10214] == 10214 && 
b[10215] == 10215 && 
b[10216] == 10216 && 
b[10217] == 10217 && 
b[10218] == 10218 && 
b[10219] == 10219 && 
b[10220] == 10220 && 
b[10221] == 10221 && 
b[10222] == 10222 && 
b[10223] == 10223 && 
b[10224] == 10224 && 
b[10225] == 10225 && 
b[10226] == 10226 && 
b[10227] == 10227 && 
b[10228] == 10228 && 
b[10229] == 10229 && 
b[10230] == 10230 && 
b[10231] == 10231 && 
b[10232] == 10232 && 
b[10233] == 10233 && 
b[10234] == 10234 && 
b[10235] == 10235 && 
b[10236] == 10236 && 
b[10237] == 10237 && 
b[10238] == 10238 && 
b[10239] == 10239 && 
b[10240] == 10240 && 
b[10241] == 10241 && 
b[10242] == 10242 && 
b[10243] == 10243 && 
b[10244] == 10244 && 
b[10245] == 10245 && 
b[10246] == 10246 && 
b[10247] == 10247 && 
b[10248] == 10248 && 
b[10249] == 10249 && 
b[10250] == 10250 && 
b[10251] == 10251 && 
b[10252] == 10252 && 
b[10253] == 10253 && 
b[10254] == 10254 && 
b[10255] == 10255 && 
b[10256] == 10256 && 
b[10257] == 10257 && 
b[10258] == 10258 && 
b[10259] == 10259 && 
b[10260] == 10260 && 
b[10261] == 10261 && 
b[10262] == 10262 && 
b[10263] == 10263 && 
b[10264] == 10264 && 
b[10265] == 10265 && 
b[10266] == 10266 && 
b[10267] == 10267 && 
b[10268] == 10268 && 
b[10269] == 10269 && 
b[10270] == 10270 && 
b[10271] == 10271 && 
b[10272] == 10272 && 
b[10273] == 10273 && 
b[10274] == 10274 && 
b[10275] == 10275 && 
b[10276] == 10276 && 
b[10277] == 10277 && 
b[10278] == 10278 && 
b[10279] == 10279 && 
b[10280] == 10280 && 
b[10281] == 10281 && 
b[10282] == 10282 && 
b[10283] == 10283 && 
b[10284] == 10284 && 
b[10285] == 10285 && 
b[10286] == 10286 && 
b[10287] == 10287 && 
b[10288] == 10288 && 
b[10289] == 10289 && 
b[10290] == 10290 && 
b[10291] == 10291 && 
b[10292] == 10292 && 
b[10293] == 10293 && 
b[10294] == 10294 && 
b[10295] == 10295 && 
b[10296] == 10296 && 
b[10297] == 10297 && 
b[10298] == 10298 && 
b[10299] == 10299 && 
b[10300] == 10300 && 
b[10301] == 10301 && 
b[10302] == 10302 && 
b[10303] == 10303 && 
b[10304] == 10304 && 
b[10305] == 10305 && 
b[10306] == 10306 && 
b[10307] == 10307 && 
b[10308] == 10308 && 
b[10309] == 10309 && 
b[10310] == 10310 && 
b[10311] == 10311 && 
b[10312] == 10312 && 
b[10313] == 10313 && 
b[10314] == 10314 && 
b[10315] == 10315 && 
b[10316] == 10316 && 
b[10317] == 10317 && 
b[10318] == 10318 && 
b[10319] == 10319 && 
b[10320] == 10320 && 
b[10321] == 10321 && 
b[10322] == 10322 && 
b[10323] == 10323 && 
b[10324] == 10324 && 
b[10325] == 10325 && 
b[10326] == 10326 && 
b[10327] == 10327 && 
b[10328] == 10328 && 
b[10329] == 10329 && 
b[10330] == 10330 && 
b[10331] == 10331 && 
b[10332] == 10332 && 
b[10333] == 10333 && 
b[10334] == 10334 && 
b[10335] == 10335 && 
b[10336] == 10336 && 
b[10337] == 10337 && 
b[10338] == 10338 && 
b[10339] == 10339 && 
b[10340] == 10340 && 
b[10341] == 10341 && 
b[10342] == 10342 && 
b[10343] == 10343 && 
b[10344] == 10344 && 
b[10345] == 10345 && 
b[10346] == 10346 && 
b[10347] == 10347 && 
b[10348] == 10348 && 
b[10349] == 10349 && 
b[10350] == 10350 && 
b[10351] == 10351 && 
b[10352] == 10352 && 
b[10353] == 10353 && 
b[10354] == 10354 && 
b[10355] == 10355 && 
b[10356] == 10356 && 
b[10357] == 10357 && 
b[10358] == 10358 && 
b[10359] == 10359 && 
b[10360] == 10360 && 
b[10361] == 10361 && 
b[10362] == 10362 && 
b[10363] == 10363 && 
b[10364] == 10364 && 
b[10365] == 10365 && 
b[10366] == 10366 && 
b[10367] == 10367 && 
b[10368] == 10368 && 
b[10369] == 10369 && 
b[10370] == 10370 && 
b[10371] == 10371 && 
b[10372] == 10372 && 
b[10373] == 10373 && 
b[10374] == 10374 && 
b[10375] == 10375 && 
b[10376] == 10376 && 
b[10377] == 10377 && 
b[10378] == 10378 && 
b[10379] == 10379 && 
b[10380] == 10380 && 
b[10381] == 10381 && 
b[10382] == 10382 && 
b[10383] == 10383 && 
b[10384] == 10384 && 
b[10385] == 10385 && 
b[10386] == 10386 && 
b[10387] == 10387 && 
b[10388] == 10388 && 
b[10389] == 10389 && 
b[10390] == 10390 && 
b[10391] == 10391 && 
b[10392] == 10392 && 
b[10393] == 10393 && 
b[10394] == 10394 && 
b[10395] == 10395 && 
b[10396] == 10396 && 
b[10397] == 10397 && 
b[10398] == 10398 && 
b[10399] == 10399 && 
b[10400] == 10400 && 
b[10401] == 10401 && 
b[10402] == 10402 && 
b[10403] == 10403 && 
b[10404] == 10404 && 
b[10405] == 10405 && 
b[10406] == 10406 && 
b[10407] == 10407 && 
b[10408] == 10408 && 
b[10409] == 10409 && 
b[10410] == 10410 && 
b[10411] == 10411 && 
b[10412] == 10412 && 
b[10413] == 10413 && 
b[10414] == 10414 && 
b[10415] == 10415 && 
b[10416] == 10416 && 
b[10417] == 10417 && 
b[10418] == 10418 && 
b[10419] == 10419 && 
b[10420] == 10420 && 
b[10421] == 10421 && 
b[10422] == 10422 && 
b[10423] == 10423 && 
b[10424] == 10424 && 
b[10425] == 10425 && 
b[10426] == 10426 && 
b[10427] == 10427 && 
b[10428] == 10428 && 
b[10429] == 10429 && 
b[10430] == 10430 && 
b[10431] == 10431 && 
b[10432] == 10432 && 
b[10433] == 10433 && 
b[10434] == 10434 && 
b[10435] == 10435 && 
b[10436] == 10436 && 
b[10437] == 10437 && 
b[10438] == 10438 && 
b[10439] == 10439 && 
b[10440] == 10440 && 
b[10441] == 10441 && 
b[10442] == 10442 && 
b[10443] == 10443 && 
b[10444] == 10444 && 
b[10445] == 10445 && 
b[10446] == 10446 && 
b[10447] == 10447 && 
b[10448] == 10448 && 
b[10449] == 10449 && 
b[10450] == 10450 && 
b[10451] == 10451 && 
b[10452] == 10452 && 
b[10453] == 10453 && 
b[10454] == 10454 && 
b[10455] == 10455 && 
b[10456] == 10456 && 
b[10457] == 10457 && 
b[10458] == 10458 && 
b[10459] == 10459 && 
b[10460] == 10460 && 
b[10461] == 10461 && 
b[10462] == 10462 && 
b[10463] == 10463 && 
b[10464] == 10464 && 
b[10465] == 10465 && 
b[10466] == 10466 && 
b[10467] == 10467 && 
b[10468] == 10468 && 
b[10469] == 10469 && 
b[10470] == 10470 && 
b[10471] == 10471 && 
b[10472] == 10472 && 
b[10473] == 10473 && 
b[10474] == 10474 && 
b[10475] == 10475 && 
b[10476] == 10476 && 
b[10477] == 10477 && 
b[10478] == 10478 && 
b[10479] == 10479 && 
b[10480] == 10480 && 
b[10481] == 10481 && 
b[10482] == 10482 && 
b[10483] == 10483 && 
b[10484] == 10484 && 
b[10485] == 10485 && 
b[10486] == 10486 && 
b[10487] == 10487 && 
b[10488] == 10488 && 
b[10489] == 10489 && 
b[10490] == 10490 && 
b[10491] == 10491 && 
b[10492] == 10492 && 
b[10493] == 10493 && 
b[10494] == 10494 && 
b[10495] == 10495 && 
b[10496] == 10496 && 
b[10497] == 10497 && 
b[10498] == 10498 && 
b[10499] == 10499 && 
b[10500] == 10500 && 
b[10501] == 10501 && 
b[10502] == 10502 && 
b[10503] == 10503 && 
b[10504] == 10504 && 
b[10505] == 10505 && 
b[10506] == 10506 && 
b[10507] == 10507 && 
b[10508] == 10508 && 
b[10509] == 10509 && 
b[10510] == 10510 && 
b[10511] == 10511 && 
b[10512] == 10512 && 
b[10513] == 10513 && 
b[10514] == 10514 && 
b[10515] == 10515 && 
b[10516] == 10516 && 
b[10517] == 10517 && 
b[10518] == 10518 && 
b[10519] == 10519 && 
b[10520] == 10520 && 
b[10521] == 10521 && 
b[10522] == 10522 && 
b[10523] == 10523 && 
b[10524] == 10524 && 
b[10525] == 10525 && 
b[10526] == 10526 && 
b[10527] == 10527 && 
b[10528] == 10528 && 
b[10529] == 10529 && 
b[10530] == 10530 && 
b[10531] == 10531 && 
b[10532] == 10532 && 
b[10533] == 10533 && 
b[10534] == 10534 && 
b[10535] == 10535 && 
b[10536] == 10536 && 
b[10537] == 10537 && 
b[10538] == 10538 && 
b[10539] == 10539 && 
b[10540] == 10540 && 
b[10541] == 10541 && 
b[10542] == 10542 && 
b[10543] == 10543 && 
b[10544] == 10544 && 
b[10545] == 10545 && 
b[10546] == 10546 && 
b[10547] == 10547 && 
b[10548] == 10548 && 
b[10549] == 10549 && 
b[10550] == 10550 && 
b[10551] == 10551 && 
b[10552] == 10552 && 
b[10553] == 10553 && 
b[10554] == 10554 && 
b[10555] == 10555 && 
b[10556] == 10556 && 
b[10557] == 10557 && 
b[10558] == 10558 && 
b[10559] == 10559 && 
b[10560] == 10560 && 
b[10561] == 10561 && 
b[10562] == 10562 && 
b[10563] == 10563 && 
b[10564] == 10564 && 
b[10565] == 10565 && 
b[10566] == 10566 && 
b[10567] == 10567 && 
b[10568] == 10568 && 
b[10569] == 10569 && 
b[10570] == 10570 && 
b[10571] == 10571 && 
b[10572] == 10572 && 
b[10573] == 10573 && 
b[10574] == 10574 && 
b[10575] == 10575 && 
b[10576] == 10576 && 
b[10577] == 10577 && 
b[10578] == 10578 && 
b[10579] == 10579 && 
b[10580] == 10580 && 
b[10581] == 10581 && 
b[10582] == 10582 && 
b[10583] == 10583 && 
b[10584] == 10584 && 
b[10585] == 10585 && 
b[10586] == 10586 && 
b[10587] == 10587 && 
b[10588] == 10588 && 
b[10589] == 10589 && 
b[10590] == 10590 && 
b[10591] == 10591 && 
b[10592] == 10592 && 
b[10593] == 10593 && 
b[10594] == 10594 && 
b[10595] == 10595 && 
b[10596] == 10596 && 
b[10597] == 10597 && 
b[10598] == 10598 && 
b[10599] == 10599 && 
b[10600] == 10600 && 
b[10601] == 10601 && 
b[10602] == 10602 && 
b[10603] == 10603 && 
b[10604] == 10604 && 
b[10605] == 10605 && 
b[10606] == 10606 && 
b[10607] == 10607 && 
b[10608] == 10608 && 
b[10609] == 10609 && 
b[10610] == 10610 && 
b[10611] == 10611 && 
b[10612] == 10612 && 
b[10613] == 10613 && 
b[10614] == 10614 && 
b[10615] == 10615 && 
b[10616] == 10616 && 
b[10617] == 10617 && 
b[10618] == 10618 && 
b[10619] == 10619 && 
b[10620] == 10620 && 
b[10621] == 10621 && 
b[10622] == 10622 && 
b[10623] == 10623 && 
b[10624] == 10624 && 
b[10625] == 10625 && 
b[10626] == 10626 && 
b[10627] == 10627 && 
b[10628] == 10628 && 
b[10629] == 10629 && 
b[10630] == 10630 && 
b[10631] == 10631 && 
b[10632] == 10632 && 
b[10633] == 10633 && 
b[10634] == 10634 && 
b[10635] == 10635 && 
b[10636] == 10636 && 
b[10637] == 10637 && 
b[10638] == 10638 && 
b[10639] == 10639 && 
b[10640] == 10640 && 
b[10641] == 10641 && 
b[10642] == 10642 && 
b[10643] == 10643 && 
b[10644] == 10644 && 
b[10645] == 10645 && 
b[10646] == 10646 && 
b[10647] == 10647 && 
b[10648] == 10648 && 
b[10649] == 10649 && 
b[10650] == 10650 && 
b[10651] == 10651 && 
b[10652] == 10652 && 
b[10653] == 10653 && 
b[10654] == 10654 && 
b[10655] == 10655 && 
b[10656] == 10656 && 
b[10657] == 10657 && 
b[10658] == 10658 && 
b[10659] == 10659 && 
b[10660] == 10660 && 
b[10661] == 10661 && 
b[10662] == 10662 && 
b[10663] == 10663 && 
b[10664] == 10664 && 
b[10665] == 10665 && 
b[10666] == 10666 && 
b[10667] == 10667 && 
b[10668] == 10668 && 
b[10669] == 10669 && 
b[10670] == 10670 && 
b[10671] == 10671 && 
b[10672] == 10672 && 
b[10673] == 10673 && 
b[10674] == 10674 && 
b[10675] == 10675 && 
b[10676] == 10676 && 
b[10677] == 10677 && 
b[10678] == 10678 && 
b[10679] == 10679 && 
b[10680] == 10680 && 
b[10681] == 10681 && 
b[10682] == 10682 && 
b[10683] == 10683 && 
b[10684] == 10684 && 
b[10685] == 10685 && 
b[10686] == 10686 && 
b[10687] == 10687 && 
b[10688] == 10688 && 
b[10689] == 10689 && 
b[10690] == 10690 && 
b[10691] == 10691 && 
b[10692] == 10692 && 
b[10693] == 10693 && 
b[10694] == 10694 && 
b[10695] == 10695 && 
b[10696] == 10696 && 
b[10697] == 10697 && 
b[10698] == 10698 && 
b[10699] == 10699 && 
b[10700] == 10700 && 
b[10701] == 10701 && 
b[10702] == 10702 && 
b[10703] == 10703 && 
b[10704] == 10704 && 
b[10705] == 10705 && 
b[10706] == 10706 && 
b[10707] == 10707 && 
b[10708] == 10708 && 
b[10709] == 10709 && 
b[10710] == 10710 && 
b[10711] == 10711 && 
b[10712] == 10712 && 
b[10713] == 10713 && 
b[10714] == 10714 && 
b[10715] == 10715 && 
b[10716] == 10716 && 
b[10717] == 10717 && 
b[10718] == 10718 && 
b[10719] == 10719 && 
b[10720] == 10720 && 
b[10721] == 10721 && 
b[10722] == 10722 && 
b[10723] == 10723 && 
b[10724] == 10724 && 
b[10725] == 10725 && 
b[10726] == 10726 && 
b[10727] == 10727 && 
b[10728] == 10728 && 
b[10729] == 10729 && 
b[10730] == 10730 && 
b[10731] == 10731 && 
b[10732] == 10732 && 
b[10733] == 10733 && 
b[10734] == 10734 && 
b[10735] == 10735 && 
b[10736] == 10736 && 
b[10737] == 10737 && 
b[10738] == 10738 && 
b[10739] == 10739 && 
b[10740] == 10740 && 
b[10741] == 10741 && 
b[10742] == 10742 && 
b[10743] == 10743 && 
b[10744] == 10744 && 
b[10745] == 10745 && 
b[10746] == 10746 && 
b[10747] == 10747 && 
b[10748] == 10748 && 
b[10749] == 10749 && 
b[10750] == 10750 && 
b[10751] == 10751 && 
b[10752] == 10752 && 
b[10753] == 10753 && 
b[10754] == 10754 && 
b[10755] == 10755 && 
b[10756] == 10756 && 
b[10757] == 10757 && 
b[10758] == 10758 && 
b[10759] == 10759 && 
b[10760] == 10760 && 
b[10761] == 10761 && 
b[10762] == 10762 && 
b[10763] == 10763 && 
b[10764] == 10764 && 
b[10765] == 10765 && 
b[10766] == 10766 && 
b[10767] == 10767 && 
b[10768] == 10768 && 
b[10769] == 10769 && 
b[10770] == 10770 && 
b[10771] == 10771 && 
b[10772] == 10772 && 
b[10773] == 10773 && 
b[10774] == 10774 && 
b[10775] == 10775 && 
b[10776] == 10776 && 
b[10777] == 10777 && 
b[10778] == 10778 && 
b[10779] == 10779 && 
b[10780] == 10780 && 
b[10781] == 10781 && 
b[10782] == 10782 && 
b[10783] == 10783 && 
b[10784] == 10784 && 
b[10785] == 10785 && 
b[10786] == 10786 && 
b[10787] == 10787 && 
b[10788] == 10788 && 
b[10789] == 10789 && 
b[10790] == 10790 && 
b[10791] == 10791 && 
b[10792] == 10792 && 
b[10793] == 10793 && 
b[10794] == 10794 && 
b[10795] == 10795 && 
b[10796] == 10796 && 
b[10797] == 10797 && 
b[10798] == 10798 && 
b[10799] == 10799 && 
b[10800] == 10800 && 
b[10801] == 10801 && 
b[10802] == 10802 && 
b[10803] == 10803 && 
b[10804] == 10804 && 
b[10805] == 10805 && 
b[10806] == 10806 && 
b[10807] == 10807 && 
b[10808] == 10808 && 
b[10809] == 10809 && 
b[10810] == 10810 && 
b[10811] == 10811 && 
b[10812] == 10812 && 
b[10813] == 10813 && 
b[10814] == 10814 && 
b[10815] == 10815 && 
b[10816] == 10816 && 
b[10817] == 10817 && 
b[10818] == 10818 && 
b[10819] == 10819 && 
b[10820] == 10820 && 
b[10821] == 10821 && 
b[10822] == 10822 && 
b[10823] == 10823 && 
b[10824] == 10824 && 
b[10825] == 10825 && 
b[10826] == 10826 && 
b[10827] == 10827 && 
b[10828] == 10828 && 
b[10829] == 10829 && 
b[10830] == 10830 && 
b[10831] == 10831 && 
b[10832] == 10832 && 
b[10833] == 10833 && 
b[10834] == 10834 && 
b[10835] == 10835 && 
b[10836] == 10836 && 
b[10837] == 10837 && 
b[10838] == 10838 && 
b[10839] == 10839 && 
b[10840] == 10840 && 
b[10841] == 10841 && 
b[10842] == 10842 && 
b[10843] == 10843 && 
b[10844] == 10844 && 
b[10845] == 10845 && 
b[10846] == 10846 && 
b[10847] == 10847 && 
b[10848] == 10848 && 
b[10849] == 10849 && 
b[10850] == 10850 && 
b[10851] == 10851 && 
b[10852] == 10852 && 
b[10853] == 10853 && 
b[10854] == 10854 && 
b[10855] == 10855 && 
b[10856] == 10856 && 
b[10857] == 10857 && 
b[10858] == 10858 && 
b[10859] == 10859 && 
b[10860] == 10860 && 
b[10861] == 10861 && 
b[10862] == 10862 && 
b[10863] == 10863 && 
b[10864] == 10864 && 
b[10865] == 10865 && 
b[10866] == 10866 && 
b[10867] == 10867 && 
b[10868] == 10868 && 
b[10869] == 10869 && 
b[10870] == 10870 && 
b[10871] == 10871 && 
b[10872] == 10872 && 
b[10873] == 10873 && 
b[10874] == 10874 && 
b[10875] == 10875 && 
b[10876] == 10876 && 
b[10877] == 10877 && 
b[10878] == 10878 && 
b[10879] == 10879 && 
b[10880] == 10880 && 
b[10881] == 10881 && 
b[10882] == 10882 && 
b[10883] == 10883 && 
b[10884] == 10884 && 
b[10885] == 10885 && 
b[10886] == 10886 && 
b[10887] == 10887 && 
b[10888] == 10888 && 
b[10889] == 10889 && 
b[10890] == 10890 && 
b[10891] == 10891 && 
b[10892] == 10892 && 
b[10893] == 10893 && 
b[10894] == 10894 && 
b[10895] == 10895 && 
b[10896] == 10896 && 
b[10897] == 10897 && 
b[10898] == 10898 && 
b[10899] == 10899 && 
b[10900] == 10900 && 
b[10901] == 10901 && 
b[10902] == 10902 && 
b[10903] == 10903 && 
b[10904] == 10904 && 
b[10905] == 10905 && 
b[10906] == 10906 && 
b[10907] == 10907 && 
b[10908] == 10908 && 
b[10909] == 10909 && 
b[10910] == 10910 && 
b[10911] == 10911 && 
b[10912] == 10912 && 
b[10913] == 10913 && 
b[10914] == 10914 && 
b[10915] == 10915 && 
b[10916] == 10916 && 
b[10917] == 10917 && 
b[10918] == 10918 && 
b[10919] == 10919 && 
b[10920] == 10920 && 
b[10921] == 10921 && 
b[10922] == 10922 && 
b[10923] == 10923 && 
b[10924] == 10924 && 
b[10925] == 10925 && 
b[10926] == 10926 && 
b[10927] == 10927 && 
b[10928] == 10928 && 
b[10929] == 10929 && 
b[10930] == 10930 && 
b[10931] == 10931 && 
b[10932] == 10932 && 
b[10933] == 10933 && 
b[10934] == 10934 && 
b[10935] == 10935 && 
b[10936] == 10936 && 
b[10937] == 10937 && 
b[10938] == 10938 && 
b[10939] == 10939 && 
b[10940] == 10940 && 
b[10941] == 10941 && 
b[10942] == 10942 && 
b[10943] == 10943 && 
b[10944] == 10944 && 
b[10945] == 10945 && 
b[10946] == 10946 && 
b[10947] == 10947 && 
b[10948] == 10948 && 
b[10949] == 10949 && 
b[10950] == 10950 && 
b[10951] == 10951 && 
b[10952] == 10952 && 
b[10953] == 10953 && 
b[10954] == 10954 && 
b[10955] == 10955 && 
b[10956] == 10956 && 
b[10957] == 10957 && 
b[10958] == 10958 && 
b[10959] == 10959 && 
b[10960] == 10960 && 
b[10961] == 10961 && 
b[10962] == 10962 && 
b[10963] == 10963 && 
b[10964] == 10964 && 
b[10965] == 10965 && 
b[10966] == 10966 && 
b[10967] == 10967 && 
b[10968] == 10968 && 
b[10969] == 10969 && 
b[10970] == 10970 && 
b[10971] == 10971 && 
b[10972] == 10972 && 
b[10973] == 10973 && 
b[10974] == 10974 && 
b[10975] == 10975 && 
b[10976] == 10976 && 
b[10977] == 10977 && 
b[10978] == 10978 && 
b[10979] == 10979 && 
b[10980] == 10980 && 
b[10981] == 10981 && 
b[10982] == 10982 && 
b[10983] == 10983 && 
b[10984] == 10984 && 
b[10985] == 10985 && 
b[10986] == 10986 && 
b[10987] == 10987 && 
b[10988] == 10988 && 
b[10989] == 10989 && 
b[10990] == 10990 && 
b[10991] == 10991 && 
b[10992] == 10992 && 
b[10993] == 10993 && 
b[10994] == 10994 && 
b[10995] == 10995 && 
b[10996] == 10996 && 
b[10997] == 10997 && 
b[10998] == 10998 && 
b[10999] == 10999 && 
b[11000] == 11000 && 
b[11001] == 11001 && 
b[11002] == 11002 && 
b[11003] == 11003 && 
b[11004] == 11004 && 
b[11005] == 11005 && 
b[11006] == 11006 && 
b[11007] == 11007 && 
b[11008] == 11008 && 
b[11009] == 11009 && 
b[11010] == 11010 && 
b[11011] == 11011 && 
b[11012] == 11012 && 
b[11013] == 11013 && 
b[11014] == 11014 && 
b[11015] == 11015 && 
b[11016] == 11016 && 
b[11017] == 11017 && 
b[11018] == 11018 && 
b[11019] == 11019 && 
b[11020] == 11020 && 
b[11021] == 11021 && 
b[11022] == 11022 && 
b[11023] == 11023 && 
b[11024] == 11024 && 
b[11025] == 11025 && 
b[11026] == 11026 && 
b[11027] == 11027 && 
b[11028] == 11028 && 
b[11029] == 11029 && 
b[11030] == 11030 && 
b[11031] == 11031 && 
b[11032] == 11032 && 
b[11033] == 11033 && 
b[11034] == 11034 && 
b[11035] == 11035 && 
b[11036] == 11036 && 
b[11037] == 11037 && 
b[11038] == 11038 && 
b[11039] == 11039 && 
b[11040] == 11040 && 
b[11041] == 11041 && 
b[11042] == 11042 && 
b[11043] == 11043 && 
b[11044] == 11044 && 
b[11045] == 11045 && 
b[11046] == 11046 && 
b[11047] == 11047 && 
b[11048] == 11048 && 
b[11049] == 11049 && 
b[11050] == 11050 && 
b[11051] == 11051 && 
b[11052] == 11052 && 
b[11053] == 11053 && 
b[11054] == 11054 && 
b[11055] == 11055 && 
b[11056] == 11056 && 
b[11057] == 11057 && 
b[11058] == 11058 && 
b[11059] == 11059 && 
b[11060] == 11060 && 
b[11061] == 11061 && 
b[11062] == 11062 && 
b[11063] == 11063 && 
b[11064] == 11064 && 
b[11065] == 11065 && 
b[11066] == 11066 && 
b[11067] == 11067 && 
b[11068] == 11068 && 
b[11069] == 11069 && 
b[11070] == 11070 && 
b[11071] == 11071 && 
b[11072] == 11072 && 
b[11073] == 11073 && 
b[11074] == 11074 && 
b[11075] == 11075 && 
b[11076] == 11076 && 
b[11077] == 11077 && 
b[11078] == 11078 && 
b[11079] == 11079 && 
b[11080] == 11080 && 
b[11081] == 11081 && 
b[11082] == 11082 && 
b[11083] == 11083 && 
b[11084] == 11084 && 
b[11085] == 11085 && 
b[11086] == 11086 && 
b[11087] == 11087 && 
b[11088] == 11088 && 
b[11089] == 11089 && 
b[11090] == 11090 && 
b[11091] == 11091 && 
b[11092] == 11092 && 
b[11093] == 11093 && 
b[11094] == 11094 && 
b[11095] == 11095 && 
b[11096] == 11096 && 
b[11097] == 11097 && 
b[11098] == 11098 && 
b[11099] == 11099 && 
b[11100] == 11100 && 
b[11101] == 11101 && 
b[11102] == 11102 && 
b[11103] == 11103 && 
b[11104] == 11104 && 
b[11105] == 11105 && 
b[11106] == 11106 && 
b[11107] == 11107 && 
b[11108] == 11108 && 
b[11109] == 11109 && 
b[11110] == 11110 && 
b[11111] == 11111 && 
b[11112] == 11112 && 
b[11113] == 11113 && 
b[11114] == 11114 && 
b[11115] == 11115 && 
b[11116] == 11116 && 
b[11117] == 11117 && 
b[11118] == 11118 && 
b[11119] == 11119 && 
b[11120] == 11120 && 
b[11121] == 11121 && 
b[11122] == 11122 && 
b[11123] == 11123 && 
b[11124] == 11124 && 
b[11125] == 11125 && 
b[11126] == 11126 && 
b[11127] == 11127 && 
b[11128] == 11128 && 
b[11129] == 11129 && 
b[11130] == 11130 && 
b[11131] == 11131 && 
b[11132] == 11132 && 
b[11133] == 11133 && 
b[11134] == 11134 && 
b[11135] == 11135 && 
b[11136] == 11136 && 
b[11137] == 11137 && 
b[11138] == 11138 && 
b[11139] == 11139 && 
b[11140] == 11140 && 
b[11141] == 11141 && 
b[11142] == 11142 && 
b[11143] == 11143 && 
b[11144] == 11144 && 
b[11145] == 11145 && 
b[11146] == 11146 && 
b[11147] == 11147 && 
b[11148] == 11148 && 
b[11149] == 11149 && 
b[11150] == 11150 && 
b[11151] == 11151 && 
b[11152] == 11152 && 
b[11153] == 11153 && 
b[11154] == 11154 && 
b[11155] == 11155 && 
b[11156] == 11156 && 
b[11157] == 11157 && 
b[11158] == 11158 && 
b[11159] == 11159 && 
b[11160] == 11160 && 
b[11161] == 11161 && 
b[11162] == 11162 && 
b[11163] == 11163 && 
b[11164] == 11164 && 
b[11165] == 11165 && 
b[11166] == 11166 && 
b[11167] == 11167 && 
b[11168] == 11168 && 
b[11169] == 11169 && 
b[11170] == 11170 && 
b[11171] == 11171 && 
b[11172] == 11172 && 
b[11173] == 11173 && 
b[11174] == 11174 && 
b[11175] == 11175 && 
b[11176] == 11176 && 
b[11177] == 11177 && 
b[11178] == 11178 && 
b[11179] == 11179 && 
b[11180] == 11180 && 
b[11181] == 11181 && 
b[11182] == 11182 && 
b[11183] == 11183 && 
b[11184] == 11184 && 
b[11185] == 11185 && 
b[11186] == 11186 && 
b[11187] == 11187 && 
b[11188] == 11188 && 
b[11189] == 11189 && 
b[11190] == 11190 && 
b[11191] == 11191 && 
b[11192] == 11192 && 
b[11193] == 11193 && 
b[11194] == 11194 && 
b[11195] == 11195 && 
b[11196] == 11196 && 
b[11197] == 11197 && 
b[11198] == 11198 && 
b[11199] == 11199 && 
b[11200] == 11200 && 
b[11201] == 11201 && 
b[11202] == 11202 && 
b[11203] == 11203 && 
b[11204] == 11204 && 
b[11205] == 11205 && 
b[11206] == 11206 && 
b[11207] == 11207 && 
b[11208] == 11208 && 
b[11209] == 11209 && 
b[11210] == 11210 && 
b[11211] == 11211 && 
b[11212] == 11212 && 
b[11213] == 11213 && 
b[11214] == 11214 && 
b[11215] == 11215 && 
b[11216] == 11216 && 
b[11217] == 11217 && 
b[11218] == 11218 && 
b[11219] == 11219 && 
b[11220] == 11220 && 
b[11221] == 11221 && 
b[11222] == 11222 && 
b[11223] == 11223 && 
b[11224] == 11224 && 
b[11225] == 11225 && 
b[11226] == 11226 && 
b[11227] == 11227 && 
b[11228] == 11228 && 
b[11229] == 11229 && 
b[11230] == 11230 && 
b[11231] == 11231 && 
b[11232] == 11232 && 
b[11233] == 11233 && 
b[11234] == 11234 && 
b[11235] == 11235 && 
b[11236] == 11236 && 
b[11237] == 11237 && 
b[11238] == 11238 && 
b[11239] == 11239 && 
b[11240] == 11240 && 
b[11241] == 11241 && 
b[11242] == 11242 && 
b[11243] == 11243 && 
b[11244] == 11244 && 
b[11245] == 11245 && 
b[11246] == 11246 && 
b[11247] == 11247 && 
b[11248] == 11248 && 
b[11249] == 11249 && 
b[11250] == 11250 && 
b[11251] == 11251 && 
b[11252] == 11252 && 
b[11253] == 11253 && 
b[11254] == 11254 && 
b[11255] == 11255 && 
b[11256] == 11256 && 
b[11257] == 11257 && 
b[11258] == 11258 && 
b[11259] == 11259 && 
b[11260] == 11260 && 
b[11261] == 11261 && 
b[11262] == 11262 && 
b[11263] == 11263 && 
b[11264] == 11264 && 
b[11265] == 11265 && 
b[11266] == 11266 && 
b[11267] == 11267 && 
b[11268] == 11268 && 
b[11269] == 11269 && 
b[11270] == 11270 && 
b[11271] == 11271 && 
b[11272] == 11272 && 
b[11273] == 11273 && 
b[11274] == 11274 && 
b[11275] == 11275 && 
b[11276] == 11276 && 
b[11277] == 11277 && 
b[11278] == 11278 && 
b[11279] == 11279 && 
b[11280] == 11280 && 
b[11281] == 11281 && 
b[11282] == 11282 && 
b[11283] == 11283 && 
b[11284] == 11284 && 
b[11285] == 11285 && 
b[11286] == 11286 && 
b[11287] == 11287 && 
b[11288] == 11288 && 
b[11289] == 11289 && 
b[11290] == 11290 && 
b[11291] == 11291 && 
b[11292] == 11292 && 
b[11293] == 11293 && 
b[11294] == 11294 && 
b[11295] == 11295 && 
b[11296] == 11296 && 
b[11297] == 11297 && 
b[11298] == 11298 && 
b[11299] == 11299 && 
b[11300] == 11300 && 
b[11301] == 11301 && 
b[11302] == 11302 && 
b[11303] == 11303 && 
b[11304] == 11304 && 
b[11305] == 11305 && 
b[11306] == 11306 && 
b[11307] == 11307 && 
b[11308] == 11308 && 
b[11309] == 11309 && 
b[11310] == 11310 && 
b[11311] == 11311 && 
b[11312] == 11312 && 
b[11313] == 11313 && 
b[11314] == 11314 && 
b[11315] == 11315 && 
b[11316] == 11316 && 
b[11317] == 11317 && 
b[11318] == 11318 && 
b[11319] == 11319 && 
b[11320] == 11320 && 
b[11321] == 11321 && 
b[11322] == 11322 && 
b[11323] == 11323 && 
b[11324] == 11324 && 
b[11325] == 11325 && 
b[11326] == 11326 && 
b[11327] == 11327 && 
b[11328] == 11328 && 
b[11329] == 11329 && 
b[11330] == 11330 && 
b[11331] == 11331 && 
b[11332] == 11332 && 
b[11333] == 11333 && 
b[11334] == 11334 && 
b[11335] == 11335 && 
b[11336] == 11336 && 
b[11337] == 11337 && 
b[11338] == 11338 && 
b[11339] == 11339 && 
b[11340] == 11340 && 
b[11341] == 11341 && 
b[11342] == 11342 && 
b[11343] == 11343 && 
b[11344] == 11344 && 
b[11345] == 11345 && 
b[11346] == 11346 && 
b[11347] == 11347 && 
b[11348] == 11348 && 
b[11349] == 11349 && 
b[11350] == 11350 && 
b[11351] == 11351 && 
b[11352] == 11352 && 
b[11353] == 11353 && 
b[11354] == 11354 && 
b[11355] == 11355 && 
b[11356] == 11356 && 
b[11357] == 11357 && 
b[11358] == 11358 && 
b[11359] == 11359 && 
b[11360] == 11360 && 
b[11361] == 11361 && 
b[11362] == 11362 && 
b[11363] == 11363 && 
b[11364] == 11364 && 
b[11365] == 11365 && 
b[11366] == 11366 && 
b[11367] == 11367 && 
b[11368] == 11368 && 
b[11369] == 11369 && 
b[11370] == 11370 && 
b[11371] == 11371 && 
b[11372] == 11372 && 
b[11373] == 11373 && 
b[11374] == 11374 && 
b[11375] == 11375 && 
b[11376] == 11376 && 
b[11377] == 11377 && 
b[11378] == 11378 && 
b[11379] == 11379 && 
b[11380] == 11380 && 
b[11381] == 11381 && 
b[11382] == 11382 && 
b[11383] == 11383 && 
b[11384] == 11384 && 
b[11385] == 11385 && 
b[11386] == 11386 && 
b[11387] == 11387 && 
b[11388] == 11388 && 
b[11389] == 11389 && 
b[11390] == 11390 && 
b[11391] == 11391 && 
b[11392] == 11392 && 
b[11393] == 11393 && 
b[11394] == 11394 && 
b[11395] == 11395 && 
b[11396] == 11396 && 
b[11397] == 11397 && 
b[11398] == 11398 && 
b[11399] == 11399 && 
b[11400] == 11400 && 
b[11401] == 11401 && 
b[11402] == 11402 && 
b[11403] == 11403 && 
b[11404] == 11404 && 
b[11405] == 11405 && 
b[11406] == 11406 && 
b[11407] == 11407 && 
b[11408] == 11408 && 
b[11409] == 11409 && 
b[11410] == 11410 && 
b[11411] == 11411 && 
b[11412] == 11412 && 
b[11413] == 11413 && 
b[11414] == 11414 && 
b[11415] == 11415 && 
b[11416] == 11416 && 
b[11417] == 11417 && 
b[11418] == 11418 && 
b[11419] == 11419 && 
b[11420] == 11420 && 
b[11421] == 11421 && 
b[11422] == 11422 && 
b[11423] == 11423 && 
b[11424] == 11424 && 
b[11425] == 11425 && 
b[11426] == 11426 && 
b[11427] == 11427 && 
b[11428] == 11428 && 
b[11429] == 11429 && 
b[11430] == 11430 && 
b[11431] == 11431 && 
b[11432] == 11432 && 
b[11433] == 11433 && 
b[11434] == 11434 && 
b[11435] == 11435 && 
b[11436] == 11436 && 
b[11437] == 11437 && 
b[11438] == 11438 && 
b[11439] == 11439 && 
b[11440] == 11440 && 
b[11441] == 11441 && 
b[11442] == 11442 && 
b[11443] == 11443 && 
b[11444] == 11444 && 
b[11445] == 11445 && 
b[11446] == 11446 && 
b[11447] == 11447 && 
b[11448] == 11448 && 
b[11449] == 11449 && 
b[11450] == 11450 && 
b[11451] == 11451 && 
b[11452] == 11452 && 
b[11453] == 11453 && 
b[11454] == 11454 && 
b[11455] == 11455 && 
b[11456] == 11456 && 
b[11457] == 11457 && 
b[11458] == 11458 && 
b[11459] == 11459 && 
b[11460] == 11460 && 
b[11461] == 11461 && 
b[11462] == 11462 && 
b[11463] == 11463 && 
b[11464] == 11464 && 
b[11465] == 11465 && 
b[11466] == 11466 && 
b[11467] == 11467 && 
b[11468] == 11468 && 
b[11469] == 11469 && 
b[11470] == 11470 && 
b[11471] == 11471 && 
b[11472] == 11472 && 
b[11473] == 11473 && 
b[11474] == 11474 && 
b[11475] == 11475 && 
b[11476] == 11476 && 
b[11477] == 11477 && 
b[11478] == 11478 && 
b[11479] == 11479 && 
b[11480] == 11480 && 
b[11481] == 11481 && 
b[11482] == 11482 && 
b[11483] == 11483 && 
b[11484] == 11484 && 
b[11485] == 11485 && 
b[11486] == 11486 && 
b[11487] == 11487 && 
b[11488] == 11488 && 
b[11489] == 11489 && 
b[11490] == 11490 && 
b[11491] == 11491 && 
b[11492] == 11492 && 
b[11493] == 11493 && 
b[11494] == 11494 && 
b[11495] == 11495 && 
b[11496] == 11496 && 
b[11497] == 11497 && 
b[11498] == 11498 && 
b[11499] == 11499 && 
b[11500] == 11500 && 
b[11501] == 11501 && 
b[11502] == 11502 && 
b[11503] == 11503 && 
b[11504] == 11504 && 
b[11505] == 11505 && 
b[11506] == 11506 && 
b[11507] == 11507 && 
b[11508] == 11508 && 
b[11509] == 11509 && 
b[11510] == 11510 && 
b[11511] == 11511 && 
b[11512] == 11512 && 
b[11513] == 11513 && 
b[11514] == 11514 && 
b[11515] == 11515 && 
b[11516] == 11516 && 
b[11517] == 11517 && 
b[11518] == 11518 && 
b[11519] == 11519 && 
b[11520] == 11520 && 
b[11521] == 11521 && 
b[11522] == 11522 && 
b[11523] == 11523 && 
b[11524] == 11524 && 
b[11525] == 11525 && 
b[11526] == 11526 && 
b[11527] == 11527 && 
b[11528] == 11528 && 
b[11529] == 11529 && 
b[11530] == 11530 && 
b[11531] == 11531 && 
b[11532] == 11532 && 
b[11533] == 11533 && 
b[11534] == 11534 && 
b[11535] == 11535 && 
b[11536] == 11536 && 
b[11537] == 11537 && 
b[11538] == 11538 && 
b[11539] == 11539 && 
b[11540] == 11540 && 
b[11541] == 11541 && 
b[11542] == 11542 && 
b[11543] == 11543 && 
b[11544] == 11544 && 
b[11545] == 11545 && 
b[11546] == 11546 && 
b[11547] == 11547 && 
b[11548] == 11548 && 
b[11549] == 11549 && 
b[11550] == 11550 && 
b[11551] == 11551 && 
b[11552] == 11552 && 
b[11553] == 11553 && 
b[11554] == 11554 && 
b[11555] == 11555 && 
b[11556] == 11556 && 
b[11557] == 11557 && 
b[11558] == 11558 && 
b[11559] == 11559 && 
b[11560] == 11560 && 
b[11561] == 11561 && 
b[11562] == 11562 && 
b[11563] == 11563 && 
b[11564] == 11564 && 
b[11565] == 11565 && 
b[11566] == 11566 && 
b[11567] == 11567 && 
b[11568] == 11568 && 
b[11569] == 11569 && 
b[11570] == 11570 && 
b[11571] == 11571 && 
b[11572] == 11572 && 
b[11573] == 11573 && 
b[11574] == 11574 && 
b[11575] == 11575 && 
b[11576] == 11576 && 
b[11577] == 11577 && 
b[11578] == 11578 && 
b[11579] == 11579 && 
b[11580] == 11580 && 
b[11581] == 11581 && 
b[11582] == 11582 && 
b[11583] == 11583 && 
b[11584] == 11584 && 
b[11585] == 11585 && 
b[11586] == 11586 && 
b[11587] == 11587 && 
b[11588] == 11588 && 
b[11589] == 11589 && 
b[11590] == 11590 && 
b[11591] == 11591 && 
b[11592] == 11592 && 
b[11593] == 11593 && 
b[11594] == 11594 && 
b[11595] == 11595 && 
b[11596] == 11596 && 
b[11597] == 11597 && 
b[11598] == 11598 && 
b[11599] == 11599 && 
b[11600] == 11600 && 
b[11601] == 11601 && 
b[11602] == 11602 && 
b[11603] == 11603 && 
b[11604] == 11604 && 
b[11605] == 11605 && 
b[11606] == 11606 && 
b[11607] == 11607 && 
b[11608] == 11608 && 
b[11609] == 11609 && 
b[11610] == 11610 && 
b[11611] == 11611 && 
b[11612] == 11612 && 
b[11613] == 11613 && 
b[11614] == 11614 && 
b[11615] == 11615 && 
b[11616] == 11616 && 
b[11617] == 11617 && 
b[11618] == 11618 && 
b[11619] == 11619 && 
b[11620] == 11620 && 
b[11621] == 11621 && 
b[11622] == 11622 && 
b[11623] == 11623 && 
b[11624] == 11624 && 
b[11625] == 11625 && 
b[11626] == 11626 && 
b[11627] == 11627 && 
b[11628] == 11628 && 
b[11629] == 11629 && 
b[11630] == 11630 && 
b[11631] == 11631 && 
b[11632] == 11632 && 
b[11633] == 11633 && 
b[11634] == 11634 && 
b[11635] == 11635 && 
b[11636] == 11636 && 
b[11637] == 11637 && 
b[11638] == 11638 && 
b[11639] == 11639 && 
b[11640] == 11640 && 
b[11641] == 11641 && 
b[11642] == 11642 && 
b[11643] == 11643 && 
b[11644] == 11644 && 
b[11645] == 11645 && 
b[11646] == 11646 && 
b[11647] == 11647 && 
b[11648] == 11648 && 
b[11649] == 11649 && 
b[11650] == 11650 && 
b[11651] == 11651 && 
b[11652] == 11652 && 
b[11653] == 11653 && 
b[11654] == 11654 && 
b[11655] == 11655 && 
b[11656] == 11656 && 
b[11657] == 11657 && 
b[11658] == 11658 && 
b[11659] == 11659 && 
b[11660] == 11660 && 
b[11661] == 11661 && 
b[11662] == 11662 && 
b[11663] == 11663 && 
b[11664] == 11664 && 
b[11665] == 11665 && 
b[11666] == 11666 && 
b[11667] == 11667 && 
b[11668] == 11668 && 
b[11669] == 11669 && 
b[11670] == 11670 && 
b[11671] == 11671 && 
b[11672] == 11672 && 
b[11673] == 11673 && 
b[11674] == 11674 && 
b[11675] == 11675 && 
b[11676] == 11676 && 
b[11677] == 11677 && 
b[11678] == 11678 && 
b[11679] == 11679 && 
b[11680] == 11680 && 
b[11681] == 11681 && 
b[11682] == 11682 && 
b[11683] == 11683 && 
b[11684] == 11684 && 
b[11685] == 11685 && 
b[11686] == 11686 && 
b[11687] == 11687 && 
b[11688] == 11688 && 
b[11689] == 11689 && 
b[11690] == 11690 && 
b[11691] == 11691 && 
b[11692] == 11692 && 
b[11693] == 11693 && 
b[11694] == 11694 && 
b[11695] == 11695 && 
b[11696] == 11696 && 
b[11697] == 11697 && 
b[11698] == 11698 && 
b[11699] == 11699 && 
b[11700] == 11700 && 
b[11701] == 11701 && 
b[11702] == 11702 && 
b[11703] == 11703 && 
b[11704] == 11704 && 
b[11705] == 11705 && 
b[11706] == 11706 && 
b[11707] == 11707 && 
b[11708] == 11708 && 
b[11709] == 11709 && 
b[11710] == 11710 && 
b[11711] == 11711 && 
b[11712] == 11712 && 
b[11713] == 11713 && 
b[11714] == 11714 && 
b[11715] == 11715 && 
b[11716] == 11716 && 
b[11717] == 11717 && 
b[11718] == 11718 && 
b[11719] == 11719 && 
b[11720] == 11720 && 
b[11721] == 11721 && 
b[11722] == 11722 && 
b[11723] == 11723 && 
b[11724] == 11724 && 
b[11725] == 11725 && 
b[11726] == 11726 && 
b[11727] == 11727 && 
b[11728] == 11728 && 
b[11729] == 11729 && 
b[11730] == 11730 && 
b[11731] == 11731 && 
b[11732] == 11732 && 
b[11733] == 11733 && 
b[11734] == 11734 && 
b[11735] == 11735 && 
b[11736] == 11736 && 
b[11737] == 11737 && 
b[11738] == 11738 && 
b[11739] == 11739 && 
b[11740] == 11740 && 
b[11741] == 11741 && 
b[11742] == 11742 && 
b[11743] == 11743 && 
b[11744] == 11744 && 
b[11745] == 11745 && 
b[11746] == 11746 && 
b[11747] == 11747 && 
b[11748] == 11748 && 
b[11749] == 11749 && 
b[11750] == 11750 && 
b[11751] == 11751 && 
b[11752] == 11752 && 
b[11753] == 11753 && 
b[11754] == 11754 && 
b[11755] == 11755 && 
b[11756] == 11756 && 
b[11757] == 11757 && 
b[11758] == 11758 && 
b[11759] == 11759 && 
b[11760] == 11760 && 
b[11761] == 11761 && 
b[11762] == 11762 && 
b[11763] == 11763 && 
b[11764] == 11764 && 
b[11765] == 11765 && 
b[11766] == 11766 && 
b[11767] == 11767 && 
b[11768] == 11768 && 
b[11769] == 11769 && 
b[11770] == 11770 && 
b[11771] == 11771 && 
b[11772] == 11772 && 
b[11773] == 11773 && 
b[11774] == 11774 && 
b[11775] == 11775 && 
b[11776] == 11776 && 
b[11777] == 11777 && 
b[11778] == 11778 && 
b[11779] == 11779 && 
b[11780] == 11780 && 
b[11781] == 11781 && 
b[11782] == 11782 && 
b[11783] == 11783 && 
b[11784] == 11784 && 
b[11785] == 11785 && 
b[11786] == 11786 && 
b[11787] == 11787 && 
b[11788] == 11788 && 
b[11789] == 11789 && 
b[11790] == 11790 && 
b[11791] == 11791 && 
b[11792] == 11792 && 
b[11793] == 11793 && 
b[11794] == 11794 && 
b[11795] == 11795 && 
b[11796] == 11796 && 
b[11797] == 11797 && 
b[11798] == 11798 && 
b[11799] == 11799 && 
b[11800] == 11800 && 
b[11801] == 11801 && 
b[11802] == 11802 && 
b[11803] == 11803 && 
b[11804] == 11804 && 
b[11805] == 11805 && 
b[11806] == 11806 && 
b[11807] == 11807 && 
b[11808] == 11808 && 
b[11809] == 11809 && 
b[11810] == 11810 && 
b[11811] == 11811 && 
b[11812] == 11812 && 
b[11813] == 11813 && 
b[11814] == 11814 && 
b[11815] == 11815 && 
b[11816] == 11816 && 
b[11817] == 11817 && 
b[11818] == 11818 && 
b[11819] == 11819 && 
b[11820] == 11820 && 
b[11821] == 11821 && 
b[11822] == 11822 && 
b[11823] == 11823 && 
b[11824] == 11824 && 
b[11825] == 11825 && 
b[11826] == 11826 && 
b[11827] == 11827 && 
b[11828] == 11828 && 
b[11829] == 11829 && 
b[11830] == 11830 && 
b[11831] == 11831 && 
b[11832] == 11832 && 
b[11833] == 11833 && 
b[11834] == 11834 && 
b[11835] == 11835 && 
b[11836] == 11836 && 
b[11837] == 11837 && 
b[11838] == 11838 && 
b[11839] == 11839 && 
b[11840] == 11840 && 
b[11841] == 11841 && 
b[11842] == 11842 && 
b[11843] == 11843 && 
b[11844] == 11844 && 
b[11845] == 11845 && 
b[11846] == 11846 && 
b[11847] == 11847 && 
b[11848] == 11848 && 
b[11849] == 11849 && 
b[11850] == 11850 && 
b[11851] == 11851 && 
b[11852] == 11852 && 
b[11853] == 11853 && 
b[11854] == 11854 && 
b[11855] == 11855 && 
b[11856] == 11856 && 
b[11857] == 11857 && 
b[11858] == 11858 && 
b[11859] == 11859 && 
b[11860] == 11860 && 
b[11861] == 11861 && 
b[11862] == 11862 && 
b[11863] == 11863 && 
b[11864] == 11864 && 
b[11865] == 11865 && 
b[11866] == 11866 && 
b[11867] == 11867 && 
b[11868] == 11868 && 
b[11869] == 11869 && 
b[11870] == 11870 && 
b[11871] == 11871 && 
b[11872] == 11872 && 
b[11873] == 11873 && 
b[11874] == 11874 && 
b[11875] == 11875 && 
b[11876] == 11876 && 
b[11877] == 11877 && 
b[11878] == 11878 && 
b[11879] == 11879 && 
b[11880] == 11880 && 
b[11881] == 11881 && 
b[11882] == 11882 && 
b[11883] == 11883 && 
b[11884] == 11884 && 
b[11885] == 11885 && 
b[11886] == 11886 && 
b[11887] == 11887 && 
b[11888] == 11888 && 
b[11889] == 11889 && 
b[11890] == 11890 && 
b[11891] == 11891 && 
b[11892] == 11892 && 
b[11893] == 11893 && 
b[11894] == 11894 && 
b[11895] == 11895 && 
b[11896] == 11896 && 
b[11897] == 11897 && 
b[11898] == 11898 && 
b[11899] == 11899 && 
b[11900] == 11900 && 
b[11901] == 11901 && 
b[11902] == 11902 && 
b[11903] == 11903 && 
b[11904] == 11904 && 
b[11905] == 11905 && 
b[11906] == 11906 && 
b[11907] == 11907 && 
b[11908] == 11908 && 
b[11909] == 11909 && 
b[11910] == 11910 && 
b[11911] == 11911 && 
b[11912] == 11912 && 
b[11913] == 11913 && 
b[11914] == 11914 && 
b[11915] == 11915 && 
b[11916] == 11916 && 
b[11917] == 11917 && 
b[11918] == 11918 && 
b[11919] == 11919 && 
b[11920] == 11920 && 
b[11921] == 11921 && 
b[11922] == 11922 && 
b[11923] == 11923 && 
b[11924] == 11924 && 
b[11925] == 11925 && 
b[11926] == 11926 && 
b[11927] == 11927 && 
b[11928] == 11928 && 
b[11929] == 11929 && 
b[11930] == 11930 && 
b[11931] == 11931 && 
b[11932] == 11932 && 
b[11933] == 11933 && 
b[11934] == 11934 && 
b[11935] == 11935 && 
b[11936] == 11936 && 
b[11937] == 11937 && 
b[11938] == 11938 && 
b[11939] == 11939 && 
b[11940] == 11940 && 
b[11941] == 11941 && 
b[11942] == 11942 && 
b[11943] == 11943 && 
b[11944] == 11944 && 
b[11945] == 11945 && 
b[11946] == 11946 && 
b[11947] == 11947 && 
b[11948] == 11948 && 
b[11949] == 11949 && 
b[11950] == 11950 && 
b[11951] == 11951 && 
b[11952] == 11952 && 
b[11953] == 11953 && 
b[11954] == 11954 && 
b[11955] == 11955 && 
b[11956] == 11956 && 
b[11957] == 11957 && 
b[11958] == 11958 && 
b[11959] == 11959 && 
b[11960] == 11960 && 
b[11961] == 11961 && 
b[11962] == 11962 && 
b[11963] == 11963 && 
b[11964] == 11964 && 
b[11965] == 11965 && 
b[11966] == 11966 && 
b[11967] == 11967 && 
b[11968] == 11968 && 
b[11969] == 11969 && 
b[11970] == 11970 && 
b[11971] == 11971 && 
b[11972] == 11972 && 
b[11973] == 11973 && 
b[11974] == 11974 && 
b[11975] == 11975 && 
b[11976] == 11976 && 
b[11977] == 11977 && 
b[11978] == 11978 && 
b[11979] == 11979 && 
b[11980] == 11980 && 
b[11981] == 11981 && 
b[11982] == 11982 && 
b[11983] == 11983 && 
b[11984] == 11984 && 
b[11985] == 11985 && 
b[11986] == 11986 && 
b[11987] == 11987 && 
b[11988] == 11988 && 
b[11989] == 11989 && 
b[11990] == 11990 && 
b[11991] == 11991 && 
b[11992] == 11992 && 
b[11993] == 11993 && 
b[11994] == 11994 && 
b[11995] == 11995 && 
b[11996] == 11996 && 
b[11997] == 11997 && 
b[11998] == 11998 && 
b[11999] == 11999 && 
b[12000] == 12000 && 
b[12001] == 12001 && 
b[12002] == 12002 && 
b[12003] == 12003 && 
b[12004] == 12004 && 
b[12005] == 12005 && 
b[12006] == 12006 && 
b[12007] == 12007 && 
b[12008] == 12008 && 
b[12009] == 12009 && 
b[12010] == 12010 && 
b[12011] == 12011 && 
b[12012] == 12012 && 
b[12013] == 12013 && 
b[12014] == 12014 && 
b[12015] == 12015 && 
b[12016] == 12016 && 
b[12017] == 12017 && 
b[12018] == 12018 && 
b[12019] == 12019 && 
b[12020] == 12020 && 
b[12021] == 12021 && 
b[12022] == 12022 && 
b[12023] == 12023 && 
b[12024] == 12024 && 
b[12025] == 12025 && 
b[12026] == 12026 && 
b[12027] == 12027 && 
b[12028] == 12028 && 
b[12029] == 12029 && 
b[12030] == 12030 && 
b[12031] == 12031 && 
b[12032] == 12032 && 
b[12033] == 12033 && 
b[12034] == 12034 && 
b[12035] == 12035 && 
b[12036] == 12036 && 
b[12037] == 12037 && 
b[12038] == 12038 && 
b[12039] == 12039 && 
b[12040] == 12040 && 
b[12041] == 12041 && 
b[12042] == 12042 && 
b[12043] == 12043 && 
b[12044] == 12044 && 
b[12045] == 12045 && 
b[12046] == 12046 && 
b[12047] == 12047 && 
b[12048] == 12048 && 
b[12049] == 12049 && 
b[12050] == 12050 && 
b[12051] == 12051 && 
b[12052] == 12052 && 
b[12053] == 12053 && 
b[12054] == 12054 && 
b[12055] == 12055 && 
b[12056] == 12056 && 
b[12057] == 12057 && 
b[12058] == 12058 && 
b[12059] == 12059 && 
b[12060] == 12060 && 
b[12061] == 12061 && 
b[12062] == 12062 && 
b[12063] == 12063 && 
b[12064] == 12064 && 
b[12065] == 12065 && 
b[12066] == 12066 && 
b[12067] == 12067 && 
b[12068] == 12068 && 
b[12069] == 12069 && 
b[12070] == 12070 && 
b[12071] == 12071 && 
b[12072] == 12072 && 
b[12073] == 12073 && 
b[12074] == 12074 && 
b[12075] == 12075 && 
b[12076] == 12076 && 
b[12077] == 12077 && 
b[12078] == 12078 && 
b[12079] == 12079 && 
b[12080] == 12080 && 
b[12081] == 12081 && 
b[12082] == 12082 && 
b[12083] == 12083 && 
b[12084] == 12084 && 
b[12085] == 12085 && 
b[12086] == 12086 && 
b[12087] == 12087 && 
b[12088] == 12088 && 
b[12089] == 12089 && 
b[12090] == 12090 && 
b[12091] == 12091 && 
b[12092] == 12092 && 
b[12093] == 12093 && 
b[12094] == 12094 && 
b[12095] == 12095 && 
b[12096] == 12096 && 
b[12097] == 12097 && 
b[12098] == 12098 && 
b[12099] == 12099 && 
b[12100] == 12100 && 
b[12101] == 12101 && 
b[12102] == 12102 && 
b[12103] == 12103 && 
b[12104] == 12104 && 
b[12105] == 12105 && 
b[12106] == 12106 && 
b[12107] == 12107 && 
b[12108] == 12108 && 
b[12109] == 12109 && 
b[12110] == 12110 && 
b[12111] == 12111 && 
b[12112] == 12112 && 
b[12113] == 12113 && 
b[12114] == 12114 && 
b[12115] == 12115 && 
b[12116] == 12116 && 
b[12117] == 12117 && 
b[12118] == 12118 && 
b[12119] == 12119 && 
b[12120] == 12120 && 
b[12121] == 12121 && 
b[12122] == 12122 && 
b[12123] == 12123 && 
b[12124] == 12124 && 
b[12125] == 12125 && 
b[12126] == 12126 && 
b[12127] == 12127 && 
b[12128] == 12128 && 
b[12129] == 12129 && 
b[12130] == 12130 && 
b[12131] == 12131 && 
b[12132] == 12132 && 
b[12133] == 12133 && 
b[12134] == 12134 && 
b[12135] == 12135 && 
b[12136] == 12136 && 
b[12137] == 12137 && 
b[12138] == 12138 && 
b[12139] == 12139 && 
b[12140] == 12140 && 
b[12141] == 12141 && 
b[12142] == 12142 && 
b[12143] == 12143 && 
b[12144] == 12144 && 
b[12145] == 12145 && 
b[12146] == 12146 && 
b[12147] == 12147 && 
b[12148] == 12148 && 
b[12149] == 12149 && 
b[12150] == 12150 && 
b[12151] == 12151 && 
b[12152] == 12152 && 
b[12153] == 12153 && 
b[12154] == 12154 && 
b[12155] == 12155 && 
b[12156] == 12156 && 
b[12157] == 12157 && 
b[12158] == 12158 && 
b[12159] == 12159 && 
b[12160] == 12160 && 
b[12161] == 12161 && 
b[12162] == 12162 && 
b[12163] == 12163 && 
b[12164] == 12164 && 
b[12165] == 12165 && 
b[12166] == 12166 && 
b[12167] == 12167 && 
b[12168] == 12168 && 
b[12169] == 12169 && 
b[12170] == 12170 && 
b[12171] == 12171 && 
b[12172] == 12172 && 
b[12173] == 12173 && 
b[12174] == 12174 && 
b[12175] == 12175 && 
b[12176] == 12176 && 
b[12177] == 12177 && 
b[12178] == 12178 && 
b[12179] == 12179 && 
b[12180] == 12180 && 
b[12181] == 12181 && 
b[12182] == 12182 && 
b[12183] == 12183 && 
b[12184] == 12184 && 
b[12185] == 12185 && 
b[12186] == 12186 && 
b[12187] == 12187 && 
b[12188] == 12188 && 
b[12189] == 12189 && 
b[12190] == 12190 && 
b[12191] == 12191 && 
b[12192] == 12192 && 
b[12193] == 12193 && 
b[12194] == 12194 && 
b[12195] == 12195 && 
b[12196] == 12196 && 
b[12197] == 12197 && 
b[12198] == 12198 && 
b[12199] == 12199 && 
b[12200] == 12200 && 
b[12201] == 12201 && 
b[12202] == 12202 && 
b[12203] == 12203 && 
b[12204] == 12204 && 
b[12205] == 12205 && 
b[12206] == 12206 && 
b[12207] == 12207 && 
b[12208] == 12208 && 
b[12209] == 12209 && 
b[12210] == 12210 && 
b[12211] == 12211 && 
b[12212] == 12212 && 
b[12213] == 12213 && 
b[12214] == 12214 && 
b[12215] == 12215 && 
b[12216] == 12216 && 
b[12217] == 12217 && 
b[12218] == 12218 && 
b[12219] == 12219 && 
b[12220] == 12220 && 
b[12221] == 12221 && 
b[12222] == 12222 && 
b[12223] == 12223 && 
b[12224] == 12224 && 
b[12225] == 12225 && 
b[12226] == 12226 && 
b[12227] == 12227 && 
b[12228] == 12228 && 
b[12229] == 12229 && 
b[12230] == 12230 && 
b[12231] == 12231 && 
b[12232] == 12232 && 
b[12233] == 12233 && 
b[12234] == 12234 && 
b[12235] == 12235 && 
b[12236] == 12236 && 
b[12237] == 12237 && 
b[12238] == 12238 && 
b[12239] == 12239 && 
b[12240] == 12240 && 
b[12241] == 12241 && 
b[12242] == 12242 && 
b[12243] == 12243 && 
b[12244] == 12244 && 
b[12245] == 12245 && 
b[12246] == 12246 && 
b[12247] == 12247 && 
b[12248] == 12248 && 
b[12249] == 12249 && 
b[12250] == 12250 && 
b[12251] == 12251 && 
b[12252] == 12252 && 
b[12253] == 12253 && 
b[12254] == 12254 && 
b[12255] == 12255 && 
b[12256] == 12256 && 
b[12257] == 12257 && 
b[12258] == 12258 && 
b[12259] == 12259 && 
b[12260] == 12260 && 
b[12261] == 12261 && 
b[12262] == 12262 && 
b[12263] == 12263 && 
b[12264] == 12264 && 
b[12265] == 12265 && 
b[12266] == 12266 && 
b[12267] == 12267 && 
b[12268] == 12268 && 
b[12269] == 12269 && 
b[12270] == 12270 && 
b[12271] == 12271 && 
b[12272] == 12272 && 
b[12273] == 12273 && 
b[12274] == 12274 && 
b[12275] == 12275 && 
b[12276] == 12276 && 
b[12277] == 12277 && 
b[12278] == 12278 && 
b[12279] == 12279 && 
b[12280] == 12280 && 
b[12281] == 12281 && 
b[12282] == 12282 && 
b[12283] == 12283 && 
b[12284] == 12284 && 
b[12285] == 12285 && 
b[12286] == 12286 && 
b[12287] == 12287 && 
b[12288] == 12288 && 
b[12289] == 12289 && 
b[12290] == 12290 && 
b[12291] == 12291 && 
b[12292] == 12292 && 
b[12293] == 12293 && 
b[12294] == 12294 && 
b[12295] == 12295 && 
b[12296] == 12296 && 
b[12297] == 12297 && 
b[12298] == 12298 && 
b[12299] == 12299 && 
b[12300] == 12300 && 
b[12301] == 12301 && 
b[12302] == 12302 && 
b[12303] == 12303 && 
b[12304] == 12304 && 
b[12305] == 12305 && 
b[12306] == 12306 && 
b[12307] == 12307 && 
b[12308] == 12308 && 
b[12309] == 12309 && 
b[12310] == 12310 && 
b[12311] == 12311 && 
b[12312] == 12312 && 
b[12313] == 12313 && 
b[12314] == 12314 && 
b[12315] == 12315 && 
b[12316] == 12316 && 
b[12317] == 12317 && 
b[12318] == 12318 && 
b[12319] == 12319 && 
b[12320] == 12320 && 
b[12321] == 12321 && 
b[12322] == 12322 && 
b[12323] == 12323 && 
b[12324] == 12324 && 
b[12325] == 12325 && 
b[12326] == 12326 && 
b[12327] == 12327 && 
b[12328] == 12328 && 
b[12329] == 12329 && 
b[12330] == 12330 && 
b[12331] == 12331 && 
b[12332] == 12332 && 
b[12333] == 12333 && 
b[12334] == 12334 && 
b[12335] == 12335 && 
b[12336] == 12336 && 
b[12337] == 12337 && 
b[12338] == 12338 && 
b[12339] == 12339 && 
b[12340] == 12340 && 
b[12341] == 12341 && 
b[12342] == 12342 && 
b[12343] == 12343 && 
b[12344] == 12344 && 
b[12345] == 12345 && 
b[12346] == 12346 && 
b[12347] == 12347 && 
b[12348] == 12348 && 
b[12349] == 12349 && 
b[12350] == 12350 && 
b[12351] == 12351 && 
b[12352] == 12352 && 
b[12353] == 12353 && 
b[12354] == 12354 && 
b[12355] == 12355 && 
b[12356] == 12356 && 
b[12357] == 12357 && 
b[12358] == 12358 && 
b[12359] == 12359 && 
b[12360] == 12360 && 
b[12361] == 12361 && 
b[12362] == 12362 && 
b[12363] == 12363 && 
b[12364] == 12364 && 
b[12365] == 12365 && 
b[12366] == 12366 && 
b[12367] == 12367 && 
b[12368] == 12368 && 
b[12369] == 12369 && 
b[12370] == 12370 && 
b[12371] == 12371 && 
b[12372] == 12372 && 
b[12373] == 12373 && 
b[12374] == 12374 && 
b[12375] == 12375 && 
b[12376] == 12376 && 
b[12377] == 12377 && 
b[12378] == 12378 && 
b[12379] == 12379 && 
b[12380] == 12380 && 
b[12381] == 12381 && 
b[12382] == 12382 && 
b[12383] == 12383 && 
b[12384] == 12384 && 
b[12385] == 12385 && 
b[12386] == 12386 && 
b[12387] == 12387 && 
b[12388] == 12388 && 
b[12389] == 12389 && 
b[12390] == 12390 && 
b[12391] == 12391 && 
b[12392] == 12392 && 
b[12393] == 12393 && 
b[12394] == 12394 && 
b[12395] == 12395 && 
b[12396] == 12396 && 
b[12397] == 12397 && 
b[12398] == 12398 && 
b[12399] == 12399 && 
b[12400] == 12400 && 
b[12401] == 12401 && 
b[12402] == 12402 && 
b[12403] == 12403 && 
b[12404] == 12404 && 
b[12405] == 12405 && 
b[12406] == 12406 && 
b[12407] == 12407 && 
b[12408] == 12408 && 
b[12409] == 12409 && 
b[12410] == 12410 && 
b[12411] == 12411 && 
b[12412] == 12412 && 
b[12413] == 12413 && 
b[12414] == 12414 && 
b[12415] == 12415 && 
b[12416] == 12416 && 
b[12417] == 12417 && 
b[12418] == 12418 && 
b[12419] == 12419 && 
b[12420] == 12420 && 
b[12421] == 12421 && 
b[12422] == 12422 && 
b[12423] == 12423 && 
b[12424] == 12424 && 
b[12425] == 12425 && 
b[12426] == 12426 && 
b[12427] == 12427 && 
b[12428] == 12428 && 
b[12429] == 12429 && 
b[12430] == 12430 && 
b[12431] == 12431 && 
b[12432] == 12432 && 
b[12433] == 12433 && 
b[12434] == 12434 && 
b[12435] == 12435 && 
b[12436] == 12436 && 
b[12437] == 12437 && 
b[12438] == 12438 && 
b[12439] == 12439 && 
b[12440] == 12440 && 
b[12441] == 12441 && 
b[12442] == 12442 && 
b[12443] == 12443 && 
b[12444] == 12444 && 
b[12445] == 12445 && 
b[12446] == 12446 && 
b[12447] == 12447 && 
b[12448] == 12448 && 
b[12449] == 12449 && 
b[12450] == 12450 && 
b[12451] == 12451 && 
b[12452] == 12452 && 
b[12453] == 12453 && 
b[12454] == 12454 && 
b[12455] == 12455 && 
b[12456] == 12456 && 
b[12457] == 12457 && 
b[12458] == 12458 && 
b[12459] == 12459 && 
b[12460] == 12460 && 
b[12461] == 12461 && 
b[12462] == 12462 && 
b[12463] == 12463 && 
b[12464] == 12464 && 
b[12465] == 12465 && 
b[12466] == 12466 && 
b[12467] == 12467 && 
b[12468] == 12468 && 
b[12469] == 12469 && 
b[12470] == 12470 && 
b[12471] == 12471 && 
b[12472] == 12472 && 
b[12473] == 12473 && 
b[12474] == 12474 && 
b[12475] == 12475 && 
b[12476] == 12476 && 
b[12477] == 12477 && 
b[12478] == 12478 && 
b[12479] == 12479 && 
b[12480] == 12480 && 
b[12481] == 12481 && 
b[12482] == 12482 && 
b[12483] == 12483 && 
b[12484] == 12484 && 
b[12485] == 12485 && 
b[12486] == 12486 && 
b[12487] == 12487 && 
b[12488] == 12488 && 
b[12489] == 12489 && 
b[12490] == 12490 && 
b[12491] == 12491 && 
b[12492] == 12492 && 
b[12493] == 12493 && 
b[12494] == 12494 && 
b[12495] == 12495 && 
b[12496] == 12496 && 
b[12497] == 12497 && 
b[12498] == 12498 && 
b[12499] == 12499 && 
b[12500] == 12500 && 
b[12501] == 12501 && 
b[12502] == 12502 && 
b[12503] == 12503 && 
b[12504] == 12504 && 
b[12505] == 12505 && 
b[12506] == 12506 && 
b[12507] == 12507 && 
b[12508] == 12508 && 
b[12509] == 12509 && 
b[12510] == 12510 && 
b[12511] == 12511 && 
b[12512] == 12512 && 
b[12513] == 12513 && 
b[12514] == 12514 && 
b[12515] == 12515 && 
b[12516] == 12516 && 
b[12517] == 12517 && 
b[12518] == 12518 && 
b[12519] == 12519 && 
b[12520] == 12520 && 
b[12521] == 12521 && 
b[12522] == 12522 && 
b[12523] == 12523 && 
b[12524] == 12524 && 
b[12525] == 12525 && 
b[12526] == 12526 && 
b[12527] == 12527 && 
b[12528] == 12528 && 
b[12529] == 12529 && 
b[12530] == 12530 && 
b[12531] == 12531 && 
b[12532] == 12532 && 
b[12533] == 12533 && 
b[12534] == 12534 && 
b[12535] == 12535 && 
b[12536] == 12536 && 
b[12537] == 12537 && 
b[12538] == 12538 && 
b[12539] == 12539 && 
b[12540] == 12540 && 
b[12541] == 12541 && 
b[12542] == 12542 && 
b[12543] == 12543 && 
b[12544] == 12544 && 
b[12545] == 12545 && 
b[12546] == 12546 && 
b[12547] == 12547 && 
b[12548] == 12548 && 
b[12549] == 12549 && 
b[12550] == 12550 && 
b[12551] == 12551 && 
b[12552] == 12552 && 
b[12553] == 12553 && 
b[12554] == 12554 && 
b[12555] == 12555 && 
b[12556] == 12556 && 
b[12557] == 12557 && 
b[12558] == 12558 && 
b[12559] == 12559 && 
b[12560] == 12560 && 
b[12561] == 12561 && 
b[12562] == 12562 && 
b[12563] == 12563 && 
b[12564] == 12564 && 
b[12565] == 12565 && 
b[12566] == 12566 && 
b[12567] == 12567 && 
b[12568] == 12568 && 
b[12569] == 12569 && 
b[12570] == 12570 && 
b[12571] == 12571 && 
b[12572] == 12572 && 
b[12573] == 12573 && 
b[12574] == 12574 && 
b[12575] == 12575 && 
b[12576] == 12576 && 
b[12577] == 12577 && 
b[12578] == 12578 && 
b[12579] == 12579 && 
b[12580] == 12580 && 
b[12581] == 12581 && 
b[12582] == 12582 && 
b[12583] == 12583 && 
b[12584] == 12584 && 
b[12585] == 12585 && 
b[12586] == 12586 && 
b[12587] == 12587 && 
b[12588] == 12588 && 
b[12589] == 12589 && 
b[12590] == 12590 && 
b[12591] == 12591 && 
b[12592] == 12592 && 
b[12593] == 12593 && 
b[12594] == 12594 && 
b[12595] == 12595 && 
b[12596] == 12596 && 
b[12597] == 12597 && 
b[12598] == 12598 && 
b[12599] == 12599 && 
b[12600] == 12600 && 
b[12601] == 12601 && 
b[12602] == 12602 && 
b[12603] == 12603 && 
b[12604] == 12604 && 
b[12605] == 12605 && 
b[12606] == 12606 && 
b[12607] == 12607 && 
b[12608] == 12608 && 
b[12609] == 12609 && 
b[12610] == 12610 && 
b[12611] == 12611 && 
b[12612] == 12612 && 
b[12613] == 12613 && 
b[12614] == 12614 && 
b[12615] == 12615 && 
b[12616] == 12616 && 
b[12617] == 12617 && 
b[12618] == 12618 && 
b[12619] == 12619 && 
b[12620] == 12620 && 
b[12621] == 12621 && 
b[12622] == 12622 && 
b[12623] == 12623 && 
b[12624] == 12624 && 
b[12625] == 12625 && 
b[12626] == 12626 && 
b[12627] == 12627 && 
b[12628] == 12628 && 
b[12629] == 12629 && 
b[12630] == 12630 && 
b[12631] == 12631 && 
b[12632] == 12632 && 
b[12633] == 12633 && 
b[12634] == 12634 && 
b[12635] == 12635 && 
b[12636] == 12636 && 
b[12637] == 12637 && 
b[12638] == 12638 && 
b[12639] == 12639 && 
b[12640] == 12640 && 
b[12641] == 12641 && 
b[12642] == 12642 && 
b[12643] == 12643 && 
b[12644] == 12644 && 
b[12645] == 12645 && 
b[12646] == 12646 && 
b[12647] == 12647 && 
b[12648] == 12648 && 
b[12649] == 12649 && 
b[12650] == 12650 && 
b[12651] == 12651 && 
b[12652] == 12652 && 
b[12653] == 12653 && 
b[12654] == 12654 && 
b[12655] == 12655 && 
b[12656] == 12656 && 
b[12657] == 12657 && 
b[12658] == 12658 && 
b[12659] == 12659 && 
b[12660] == 12660 && 
b[12661] == 12661 && 
b[12662] == 12662 && 
b[12663] == 12663 && 
b[12664] == 12664 && 
b[12665] == 12665 && 
b[12666] == 12666 && 
b[12667] == 12667 && 
b[12668] == 12668 && 
b[12669] == 12669 && 
b[12670] == 12670 && 
b[12671] == 12671 && 
b[12672] == 12672 && 
b[12673] == 12673 && 
b[12674] == 12674 && 
b[12675] == 12675 && 
b[12676] == 12676 && 
b[12677] == 12677 && 
b[12678] == 12678 && 
b[12679] == 12679 && 
b[12680] == 12680 && 
b[12681] == 12681 && 
b[12682] == 12682 && 
b[12683] == 12683 && 
b[12684] == 12684 && 
b[12685] == 12685 && 
b[12686] == 12686 && 
b[12687] == 12687 && 
b[12688] == 12688 && 
b[12689] == 12689 && 
b[12690] == 12690 && 
b[12691] == 12691 && 
b[12692] == 12692 && 
b[12693] == 12693 && 
b[12694] == 12694 && 
b[12695] == 12695 && 
b[12696] == 12696 && 
b[12697] == 12697 && 
b[12698] == 12698 && 
b[12699] == 12699 && 
b[12700] == 12700 && 
b[12701] == 12701 && 
b[12702] == 12702 && 
b[12703] == 12703 && 
b[12704] == 12704 && 
b[12705] == 12705 && 
b[12706] == 12706 && 
b[12707] == 12707 && 
b[12708] == 12708 && 
b[12709] == 12709 && 
b[12710] == 12710 && 
b[12711] == 12711 && 
b[12712] == 12712 && 
b[12713] == 12713 && 
b[12714] == 12714 && 
b[12715] == 12715 && 
b[12716] == 12716 && 
b[12717] == 12717 && 
b[12718] == 12718 && 
b[12719] == 12719 && 
b[12720] == 12720 && 
b[12721] == 12721 && 
b[12722] == 12722 && 
b[12723] == 12723 && 
b[12724] == 12724 && 
b[12725] == 12725 && 
b[12726] == 12726 && 
b[12727] == 12727 && 
b[12728] == 12728 && 
b[12729] == 12729 && 
b[12730] == 12730 && 
b[12731] == 12731 && 
b[12732] == 12732 && 
b[12733] == 12733 && 
b[12734] == 12734 && 
b[12735] == 12735 && 
b[12736] == 12736 && 
b[12737] == 12737 && 
b[12738] == 12738 && 
b[12739] == 12739 && 
b[12740] == 12740 && 
b[12741] == 12741 && 
b[12742] == 12742 && 
b[12743] == 12743 && 
b[12744] == 12744 && 
b[12745] == 12745 && 
b[12746] == 12746 && 
b[12747] == 12747 && 
b[12748] == 12748 && 
b[12749] == 12749 && 
b[12750] == 12750 && 
b[12751] == 12751 && 
b[12752] == 12752 && 
b[12753] == 12753 && 
b[12754] == 12754 && 
b[12755] == 12755 && 
b[12756] == 12756 && 
b[12757] == 12757 && 
b[12758] == 12758 && 
b[12759] == 12759 && 
b[12760] == 12760 && 
b[12761] == 12761 && 
b[12762] == 12762 && 
b[12763] == 12763 && 
b[12764] == 12764 && 
b[12765] == 12765 && 
b[12766] == 12766 && 
b[12767] == 12767 && 
b[12768] == 12768 && 
b[12769] == 12769 && 
b[12770] == 12770 && 
b[12771] == 12771 && 
b[12772] == 12772 && 
b[12773] == 12773 && 
b[12774] == 12774 && 
b[12775] == 12775 && 
b[12776] == 12776 && 
b[12777] == 12777 && 
b[12778] == 12778 && 
b[12779] == 12779 && 
b[12780] == 12780 && 
b[12781] == 12781 && 
b[12782] == 12782 && 
b[12783] == 12783 && 
b[12784] == 12784 && 
b[12785] == 12785 && 
b[12786] == 12786 && 
b[12787] == 12787 && 
b[12788] == 12788 && 
b[12789] == 12789 && 
b[12790] == 12790 && 
b[12791] == 12791 && 
b[12792] == 12792 && 
b[12793] == 12793 && 
b[12794] == 12794 && 
b[12795] == 12795 && 
b[12796] == 12796 && 
b[12797] == 12797 && 
b[12798] == 12798 && 
b[12799] == 12799 && 
b[12800] == 12800 && 
b[12801] == 12801 && 
b[12802] == 12802 && 
b[12803] == 12803 && 
b[12804] == 12804 && 
b[12805] == 12805 && 
b[12806] == 12806 && 
b[12807] == 12807 && 
b[12808] == 12808 && 
b[12809] == 12809 && 
b[12810] == 12810 && 
b[12811] == 12811 && 
b[12812] == 12812 && 
b[12813] == 12813 && 
b[12814] == 12814 && 
b[12815] == 12815 && 
b[12816] == 12816 && 
b[12817] == 12817 && 
b[12818] == 12818 && 
b[12819] == 12819 && 
b[12820] == 12820 && 
b[12821] == 12821 && 
b[12822] == 12822 && 
b[12823] == 12823 && 
b[12824] == 12824 && 
b[12825] == 12825 && 
b[12826] == 12826 && 
b[12827] == 12827 && 
b[12828] == 12828 && 
b[12829] == 12829 && 
b[12830] == 12830 && 
b[12831] == 12831 && 
b[12832] == 12832 && 
b[12833] == 12833 && 
b[12834] == 12834 && 
b[12835] == 12835 && 
b[12836] == 12836 && 
b[12837] == 12837 && 
b[12838] == 12838 && 
b[12839] == 12839 && 
b[12840] == 12840 && 
b[12841] == 12841 && 
b[12842] == 12842 && 
b[12843] == 12843 && 
b[12844] == 12844 && 
b[12845] == 12845 && 
b[12846] == 12846 && 
b[12847] == 12847 && 
b[12848] == 12848 && 
b[12849] == 12849 && 
b[12850] == 12850 && 
b[12851] == 12851 && 
b[12852] == 12852 && 
b[12853] == 12853 && 
b[12854] == 12854 && 
b[12855] == 12855 && 
b[12856] == 12856 && 
b[12857] == 12857 && 
b[12858] == 12858 && 
b[12859] == 12859 && 
b[12860] == 12860 && 
b[12861] == 12861 && 
b[12862] == 12862 && 
b[12863] == 12863 && 
b[12864] == 12864 && 
b[12865] == 12865 && 
b[12866] == 12866 && 
b[12867] == 12867 && 
b[12868] == 12868 && 
b[12869] == 12869 && 
b[12870] == 12870 && 
b[12871] == 12871 && 
b[12872] == 12872 && 
b[12873] == 12873 && 
b[12874] == 12874 && 
b[12875] == 12875 && 
b[12876] == 12876 && 
b[12877] == 12877 && 
b[12878] == 12878 && 
b[12879] == 12879 && 
b[12880] == 12880 && 
b[12881] == 12881 && 
b[12882] == 12882 && 
b[12883] == 12883 && 
b[12884] == 12884 && 
b[12885] == 12885 && 
b[12886] == 12886 && 
b[12887] == 12887 && 
b[12888] == 12888 && 
b[12889] == 12889 && 
b[12890] == 12890 && 
b[12891] == 12891 && 
b[12892] == 12892 && 
b[12893] == 12893 && 
b[12894] == 12894 && 
b[12895] == 12895 && 
b[12896] == 12896 && 
b[12897] == 12897 && 
b[12898] == 12898 && 
b[12899] == 12899 && 
b[12900] == 12900 && 
b[12901] == 12901 && 
b[12902] == 12902 && 
b[12903] == 12903 && 
b[12904] == 12904 && 
b[12905] == 12905 && 
b[12906] == 12906 && 
b[12907] == 12907 && 
b[12908] == 12908 && 
b[12909] == 12909 && 
b[12910] == 12910 && 
b[12911] == 12911 && 
b[12912] == 12912 && 
b[12913] == 12913 && 
b[12914] == 12914 && 
b[12915] == 12915 && 
b[12916] == 12916 && 
b[12917] == 12917 && 
b[12918] == 12918 && 
b[12919] == 12919 && 
b[12920] == 12920 && 
b[12921] == 12921 && 
b[12922] == 12922 && 
b[12923] == 12923 && 
b[12924] == 12924 && 
b[12925] == 12925 && 
b[12926] == 12926 && 
b[12927] == 12927 && 
b[12928] == 12928 && 
b[12929] == 12929 && 
b[12930] == 12930 && 
b[12931] == 12931 && 
b[12932] == 12932 && 
b[12933] == 12933 && 
b[12934] == 12934 && 
b[12935] == 12935 && 
b[12936] == 12936 && 
b[12937] == 12937 && 
b[12938] == 12938 && 
b[12939] == 12939 && 
b[12940] == 12940 && 
b[12941] == 12941 && 
b[12942] == 12942 && 
b[12943] == 12943 && 
b[12944] == 12944 && 
b[12945] == 12945 && 
b[12946] == 12946 && 
b[12947] == 12947 && 
b[12948] == 12948 && 
b[12949] == 12949 && 
b[12950] == 12950 && 
b[12951] == 12951 && 
b[12952] == 12952 && 
b[12953] == 12953 && 
b[12954] == 12954 && 
b[12955] == 12955 && 
b[12956] == 12956 && 
b[12957] == 12957 && 
b[12958] == 12958 && 
b[12959] == 12959 && 
b[12960] == 12960 && 
b[12961] == 12961 && 
b[12962] == 12962 && 
b[12963] == 12963 && 
b[12964] == 12964 && 
b[12965] == 12965 && 
b[12966] == 12966 && 
b[12967] == 12967 && 
b[12968] == 12968 && 
b[12969] == 12969 && 
b[12970] == 12970 && 
b[12971] == 12971 && 
b[12972] == 12972 && 
b[12973] == 12973 && 
b[12974] == 12974 && 
b[12975] == 12975 && 
b[12976] == 12976 && 
b[12977] == 12977 && 
b[12978] == 12978 && 
b[12979] == 12979 && 
b[12980] == 12980 && 
b[12981] == 12981 && 
b[12982] == 12982 && 
b[12983] == 12983 && 
b[12984] == 12984 && 
b[12985] == 12985 && 
b[12986] == 12986 && 
b[12987] == 12987 && 
b[12988] == 12988 && 
b[12989] == 12989 && 
b[12990] == 12990 && 
b[12991] == 12991 && 
b[12992] == 12992 && 
b[12993] == 12993 && 
b[12994] == 12994 && 
b[12995] == 12995 && 
b[12996] == 12996 && 
b[12997] == 12997 && 
b[12998] == 12998 && 
b[12999] == 12999 && 
b[13000] == 13000 && 
b[13001] == 13001 && 
b[13002] == 13002 && 
b[13003] == 13003 && 
b[13004] == 13004 && 
b[13005] == 13005 && 
b[13006] == 13006 && 
b[13007] == 13007 && 
b[13008] == 13008 && 
b[13009] == 13009 && 
b[13010] == 13010 && 
b[13011] == 13011 && 
b[13012] == 13012 && 
b[13013] == 13013 && 
b[13014] == 13014 && 
b[13015] == 13015 && 
b[13016] == 13016 && 
b[13017] == 13017 && 
b[13018] == 13018 && 
b[13019] == 13019 && 
b[13020] == 13020 && 
b[13021] == 13021 && 
b[13022] == 13022 && 
b[13023] == 13023 && 
b[13024] == 13024 && 
b[13025] == 13025 && 
b[13026] == 13026 && 
b[13027] == 13027 && 
b[13028] == 13028 && 
b[13029] == 13029 && 
b[13030] == 13030 && 
b[13031] == 13031 && 
b[13032] == 13032 && 
b[13033] == 13033 && 
b[13034] == 13034 && 
b[13035] == 13035 && 
b[13036] == 13036 && 
b[13037] == 13037 && 
b[13038] == 13038 && 
b[13039] == 13039 && 
b[13040] == 13040 && 
b[13041] == 13041 && 
b[13042] == 13042 && 
b[13043] == 13043 && 
b[13044] == 13044 && 
b[13045] == 13045 && 
b[13046] == 13046 && 
b[13047] == 13047 && 
b[13048] == 13048 && 
b[13049] == 13049 && 
b[13050] == 13050 && 
b[13051] == 13051 && 
b[13052] == 13052 && 
b[13053] == 13053 && 
b[13054] == 13054 && 
b[13055] == 13055 && 
b[13056] == 13056 && 
b[13057] == 13057 && 
b[13058] == 13058 && 
b[13059] == 13059 && 
b[13060] == 13060 && 
b[13061] == 13061 && 
b[13062] == 13062 && 
b[13063] == 13063 && 
b[13064] == 13064 && 
b[13065] == 13065 && 
b[13066] == 13066 && 
b[13067] == 13067 && 
b[13068] == 13068 && 
b[13069] == 13069 && 
b[13070] == 13070 && 
b[13071] == 13071 && 
b[13072] == 13072 && 
b[13073] == 13073 && 
b[13074] == 13074 && 
b[13075] == 13075 && 
b[13076] == 13076 && 
b[13077] == 13077 && 
b[13078] == 13078 && 
b[13079] == 13079 && 
b[13080] == 13080 && 
b[13081] == 13081 && 
b[13082] == 13082 && 
b[13083] == 13083 && 
b[13084] == 13084 && 
b[13085] == 13085 && 
b[13086] == 13086 && 
b[13087] == 13087 && 
b[13088] == 13088 && 
b[13089] == 13089 && 
b[13090] == 13090 && 
b[13091] == 13091 && 
b[13092] == 13092 && 
b[13093] == 13093 && 
b[13094] == 13094 && 
b[13095] == 13095 && 
b[13096] == 13096 && 
b[13097] == 13097 && 
b[13098] == 13098 && 
b[13099] == 13099 && 
b[13100] == 13100 && 
b[13101] == 13101 && 
b[13102] == 13102 && 
b[13103] == 13103 && 
b[13104] == 13104 && 
b[13105] == 13105 && 
b[13106] == 13106 && 
b[13107] == 13107 && 
b[13108] == 13108 && 
b[13109] == 13109 && 
b[13110] == 13110 && 
b[13111] == 13111 && 
b[13112] == 13112 && 
b[13113] == 13113 && 
b[13114] == 13114 && 
b[13115] == 13115 && 
b[13116] == 13116 && 
b[13117] == 13117 && 
b[13118] == 13118 && 
b[13119] == 13119 && 
b[13120] == 13120 && 
b[13121] == 13121 && 
b[13122] == 13122 && 
b[13123] == 13123 && 
b[13124] == 13124 && 
b[13125] == 13125 && 
b[13126] == 13126 && 
b[13127] == 13127 && 
b[13128] == 13128 && 
b[13129] == 13129 && 
b[13130] == 13130 && 
b[13131] == 13131 && 
b[13132] == 13132 && 
b[13133] == 13133 && 
b[13134] == 13134 && 
b[13135] == 13135 && 
b[13136] == 13136 && 
b[13137] == 13137 && 
b[13138] == 13138 && 
b[13139] == 13139 && 
b[13140] == 13140 && 
b[13141] == 13141 && 
b[13142] == 13142 && 
b[13143] == 13143 && 
b[13144] == 13144 && 
b[13145] == 13145 && 
b[13146] == 13146 && 
b[13147] == 13147 && 
b[13148] == 13148 && 
b[13149] == 13149 && 
b[13150] == 13150 && 
b[13151] == 13151 && 
b[13152] == 13152 && 
b[13153] == 13153 && 
b[13154] == 13154 && 
b[13155] == 13155 && 
b[13156] == 13156 && 
b[13157] == 13157 && 
b[13158] == 13158 && 
b[13159] == 13159 && 
b[13160] == 13160 && 
b[13161] == 13161 && 
b[13162] == 13162 && 
b[13163] == 13163 && 
b[13164] == 13164 && 
b[13165] == 13165 && 
b[13166] == 13166 && 
b[13167] == 13167 && 
b[13168] == 13168 && 
b[13169] == 13169 && 
b[13170] == 13170 && 
b[13171] == 13171 && 
b[13172] == 13172 && 
b[13173] == 13173 && 
b[13174] == 13174 && 
b[13175] == 13175 && 
b[13176] == 13176 && 
b[13177] == 13177 && 
b[13178] == 13178 && 
b[13179] == 13179 && 
b[13180] == 13180 && 
b[13181] == 13181 && 
b[13182] == 13182 && 
b[13183] == 13183 && 
b[13184] == 13184 && 
b[13185] == 13185 && 
b[13186] == 13186 && 
b[13187] == 13187 && 
b[13188] == 13188 && 
b[13189] == 13189 && 
b[13190] == 13190 && 
b[13191] == 13191 && 
b[13192] == 13192 && 
b[13193] == 13193 && 
b[13194] == 13194 && 
b[13195] == 13195 && 
b[13196] == 13196 && 
b[13197] == 13197 && 
b[13198] == 13198 && 
b[13199] == 13199 && 
b[13200] == 13200 && 
b[13201] == 13201 && 
b[13202] == 13202 && 
b[13203] == 13203 && 
b[13204] == 13204 && 
b[13205] == 13205 && 
b[13206] == 13206 && 
b[13207] == 13207 && 
b[13208] == 13208 && 
b[13209] == 13209 && 
b[13210] == 13210 && 
b[13211] == 13211 && 
b[13212] == 13212 && 
b[13213] == 13213 && 
b[13214] == 13214 && 
b[13215] == 13215 && 
b[13216] == 13216 && 
b[13217] == 13217 && 
b[13218] == 13218 && 
b[13219] == 13219 && 
b[13220] == 13220 && 
b[13221] == 13221 && 
b[13222] == 13222 && 
b[13223] == 13223 && 
b[13224] == 13224 && 
b[13225] == 13225 && 
b[13226] == 13226 && 
b[13227] == 13227 && 
b[13228] == 13228 && 
b[13229] == 13229 && 
b[13230] == 13230 && 
b[13231] == 13231 && 
b[13232] == 13232 && 
b[13233] == 13233 && 
b[13234] == 13234 && 
b[13235] == 13235 && 
b[13236] == 13236 && 
b[13237] == 13237 && 
b[13238] == 13238 && 
b[13239] == 13239 && 
b[13240] == 13240 && 
b[13241] == 13241 && 
b[13242] == 13242 && 
b[13243] == 13243 && 
b[13244] == 13244 && 
b[13245] == 13245 && 
b[13246] == 13246 && 
b[13247] == 13247 && 
b[13248] == 13248 && 
b[13249] == 13249 && 
b[13250] == 13250 && 
b[13251] == 13251 && 
b[13252] == 13252 && 
b[13253] == 13253 && 
b[13254] == 13254 && 
b[13255] == 13255 && 
b[13256] == 13256 && 
b[13257] == 13257 && 
b[13258] == 13258 && 
b[13259] == 13259 && 
b[13260] == 13260 && 
b[13261] == 13261 && 
b[13262] == 13262 && 
b[13263] == 13263 && 
b[13264] == 13264 && 
b[13265] == 13265 && 
b[13266] == 13266 && 
b[13267] == 13267 && 
b[13268] == 13268 && 
b[13269] == 13269 && 
b[13270] == 13270 && 
b[13271] == 13271 && 
b[13272] == 13272 && 
b[13273] == 13273 && 
b[13274] == 13274 && 
b[13275] == 13275 && 
b[13276] == 13276 && 
b[13277] == 13277 && 
b[13278] == 13278 && 
b[13279] == 13279 && 
b[13280] == 13280 && 
b[13281] == 13281 && 
b[13282] == 13282 && 
b[13283] == 13283 && 
b[13284] == 13284 && 
b[13285] == 13285 && 
b[13286] == 13286 && 
b[13287] == 13287 && 
b[13288] == 13288 && 
b[13289] == 13289 && 
b[13290] == 13290 && 
b[13291] == 13291 && 
b[13292] == 13292 && 
b[13293] == 13293 && 
b[13294] == 13294 && 
b[13295] == 13295 && 
b[13296] == 13296 && 
b[13297] == 13297 && 
b[13298] == 13298 && 
b[13299] == 13299 && 
b[13300] == 13300 && 
b[13301] == 13301 && 
b[13302] == 13302 && 
b[13303] == 13303 && 
b[13304] == 13304 && 
b[13305] == 13305 && 
b[13306] == 13306 && 
b[13307] == 13307 && 
b[13308] == 13308 && 
b[13309] == 13309 && 
b[13310] == 13310 && 
b[13311] == 13311 && 
b[13312] == 13312 && 
b[13313] == 13313 && 
b[13314] == 13314 && 
b[13315] == 13315 && 
b[13316] == 13316 && 
b[13317] == 13317 && 
b[13318] == 13318 && 
b[13319] == 13319 && 
b[13320] == 13320 && 
b[13321] == 13321 && 
b[13322] == 13322 && 
b[13323] == 13323 && 
b[13324] == 13324 && 
b[13325] == 13325 && 
b[13326] == 13326 && 
b[13327] == 13327 && 
b[13328] == 13328 && 
b[13329] == 13329 && 
b[13330] == 13330 && 
b[13331] == 13331 && 
b[13332] == 13332 && 
b[13333] == 13333 && 
b[13334] == 13334 && 
b[13335] == 13335 && 
b[13336] == 13336 && 
b[13337] == 13337 && 
b[13338] == 13338 && 
b[13339] == 13339 && 
b[13340] == 13340 && 
b[13341] == 13341 && 
b[13342] == 13342 && 
b[13343] == 13343 && 
b[13344] == 13344 && 
b[13345] == 13345 && 
b[13346] == 13346 && 
b[13347] == 13347 && 
b[13348] == 13348 && 
b[13349] == 13349 && 
b[13350] == 13350 && 
b[13351] == 13351 && 
b[13352] == 13352 && 
b[13353] == 13353 && 
b[13354] == 13354 && 
b[13355] == 13355 && 
b[13356] == 13356 && 
b[13357] == 13357 && 
b[13358] == 13358 && 
b[13359] == 13359 && 
b[13360] == 13360 && 
b[13361] == 13361 && 
b[13362] == 13362 && 
b[13363] == 13363 && 
b[13364] == 13364 && 
b[13365] == 13365 && 
b[13366] == 13366 && 
b[13367] == 13367 && 
b[13368] == 13368 && 
b[13369] == 13369 && 
b[13370] == 13370 && 
b[13371] == 13371 && 
b[13372] == 13372 && 
b[13373] == 13373 && 
b[13374] == 13374 && 
b[13375] == 13375 && 
b[13376] == 13376 && 
b[13377] == 13377 && 
b[13378] == 13378 && 
b[13379] == 13379 && 
b[13380] == 13380 && 
b[13381] == 13381 && 
b[13382] == 13382 && 
b[13383] == 13383 && 
b[13384] == 13384 && 
b[13385] == 13385 && 
b[13386] == 13386 && 
b[13387] == 13387 && 
b[13388] == 13388 && 
b[13389] == 13389 && 
b[13390] == 13390 && 
b[13391] == 13391 && 
b[13392] == 13392 && 
b[13393] == 13393 && 
b[13394] == 13394 && 
b[13395] == 13395 && 
b[13396] == 13396 && 
b[13397] == 13397 && 
b[13398] == 13398 && 
b[13399] == 13399 && 
b[13400] == 13400 && 
b[13401] == 13401 && 
b[13402] == 13402 && 
b[13403] == 13403 && 
b[13404] == 13404 && 
b[13405] == 13405 && 
b[13406] == 13406 && 
b[13407] == 13407 && 
b[13408] == 13408 && 
b[13409] == 13409 && 
b[13410] == 13410 && 
b[13411] == 13411 && 
b[13412] == 13412 && 
b[13413] == 13413 && 
b[13414] == 13414 && 
b[13415] == 13415 && 
b[13416] == 13416 && 
b[13417] == 13417 && 
b[13418] == 13418 && 
b[13419] == 13419 && 
b[13420] == 13420 && 
b[13421] == 13421 && 
b[13422] == 13422 && 
b[13423] == 13423 && 
b[13424] == 13424 && 
b[13425] == 13425 && 
b[13426] == 13426 && 
b[13427] == 13427 && 
b[13428] == 13428 && 
b[13429] == 13429 && 
b[13430] == 13430 && 
b[13431] == 13431 && 
b[13432] == 13432 && 
b[13433] == 13433 && 
b[13434] == 13434 && 
b[13435] == 13435 && 
b[13436] == 13436 && 
b[13437] == 13437 && 
b[13438] == 13438 && 
b[13439] == 13439 && 
b[13440] == 13440 && 
b[13441] == 13441 && 
b[13442] == 13442 && 
b[13443] == 13443 && 
b[13444] == 13444 && 
b[13445] == 13445 && 
b[13446] == 13446 && 
b[13447] == 13447 && 
b[13448] == 13448 && 
b[13449] == 13449 && 
b[13450] == 13450 && 
b[13451] == 13451 && 
b[13452] == 13452 && 
b[13453] == 13453 && 
b[13454] == 13454 && 
b[13455] == 13455 && 
b[13456] == 13456 && 
b[13457] == 13457 && 
b[13458] == 13458 && 
b[13459] == 13459 && 
b[13460] == 13460 && 
b[13461] == 13461 && 
b[13462] == 13462 && 
b[13463] == 13463 && 
b[13464] == 13464 && 
b[13465] == 13465 && 
b[13466] == 13466 && 
b[13467] == 13467 && 
b[13468] == 13468 && 
b[13469] == 13469 && 
b[13470] == 13470 && 
b[13471] == 13471 && 
b[13472] == 13472 && 
b[13473] == 13473 && 
b[13474] == 13474 && 
b[13475] == 13475 && 
b[13476] == 13476 && 
b[13477] == 13477 && 
b[13478] == 13478 && 
b[13479] == 13479 && 
b[13480] == 13480 && 
b[13481] == 13481 && 
b[13482] == 13482 && 
b[13483] == 13483 && 
b[13484] == 13484 && 
b[13485] == 13485 && 
b[13486] == 13486 && 
b[13487] == 13487 && 
b[13488] == 13488 && 
b[13489] == 13489 && 
b[13490] == 13490 && 
b[13491] == 13491 && 
b[13492] == 13492 && 
b[13493] == 13493 && 
b[13494] == 13494 && 
b[13495] == 13495 && 
b[13496] == 13496 && 
b[13497] == 13497 && 
b[13498] == 13498 && 
b[13499] == 13499 && 
b[13500] == 13500 && 
b[13501] == 13501 && 
b[13502] == 13502 && 
b[13503] == 13503 && 
b[13504] == 13504 && 
b[13505] == 13505 && 
b[13506] == 13506 && 
b[13507] == 13507 && 
b[13508] == 13508 && 
b[13509] == 13509 && 
b[13510] == 13510 && 
b[13511] == 13511 && 
b[13512] == 13512 && 
b[13513] == 13513 && 
b[13514] == 13514 && 
b[13515] == 13515 && 
b[13516] == 13516 && 
b[13517] == 13517 && 
b[13518] == 13518 && 
b[13519] == 13519 && 
b[13520] == 13520 && 
b[13521] == 13521 && 
b[13522] == 13522 && 
b[13523] == 13523 && 
b[13524] == 13524 && 
b[13525] == 13525 && 
b[13526] == 13526 && 
b[13527] == 13527 && 
b[13528] == 13528 && 
b[13529] == 13529 && 
b[13530] == 13530 && 
b[13531] == 13531 && 
b[13532] == 13532 && 
b[13533] == 13533 && 
b[13534] == 13534 && 
b[13535] == 13535 && 
b[13536] == 13536 && 
b[13537] == 13537 && 
b[13538] == 13538 && 
b[13539] == 13539 && 
b[13540] == 13540 && 
b[13541] == 13541 && 
b[13542] == 13542 && 
b[13543] == 13543 && 
b[13544] == 13544 && 
b[13545] == 13545 && 
b[13546] == 13546 && 
b[13547] == 13547 && 
b[13548] == 13548 && 
b[13549] == 13549 && 
b[13550] == 13550 && 
b[13551] == 13551 && 
b[13552] == 13552 && 
b[13553] == 13553 && 
b[13554] == 13554 && 
b[13555] == 13555 && 
b[13556] == 13556 && 
b[13557] == 13557 && 
b[13558] == 13558 && 
b[13559] == 13559 && 
b[13560] == 13560 && 
b[13561] == 13561 && 
b[13562] == 13562 && 
b[13563] == 13563 && 
b[13564] == 13564 && 
b[13565] == 13565 && 
b[13566] == 13566 && 
b[13567] == 13567 && 
b[13568] == 13568 && 
b[13569] == 13569 && 
b[13570] == 13570 && 
b[13571] == 13571 && 
b[13572] == 13572 && 
b[13573] == 13573 && 
b[13574] == 13574 && 
b[13575] == 13575 && 
b[13576] == 13576 && 
b[13577] == 13577 && 
b[13578] == 13578 && 
b[13579] == 13579 && 
b[13580] == 13580 && 
b[13581] == 13581 && 
b[13582] == 13582 && 
b[13583] == 13583 && 
b[13584] == 13584 && 
b[13585] == 13585 && 
b[13586] == 13586 && 
b[13587] == 13587 && 
b[13588] == 13588 && 
b[13589] == 13589 && 
b[13590] == 13590 && 
b[13591] == 13591 && 
b[13592] == 13592 && 
b[13593] == 13593 && 
b[13594] == 13594 && 
b[13595] == 13595 && 
b[13596] == 13596 && 
b[13597] == 13597 && 
b[13598] == 13598 && 
b[13599] == 13599 && 
b[13600] == 13600 && 
b[13601] == 13601 && 
b[13602] == 13602 && 
b[13603] == 13603 && 
b[13604] == 13604 && 
b[13605] == 13605 && 
b[13606] == 13606 && 
b[13607] == 13607 && 
b[13608] == 13608 && 
b[13609] == 13609 && 
b[13610] == 13610 && 
b[13611] == 13611 && 
b[13612] == 13612 && 
b[13613] == 13613 && 
b[13614] == 13614 && 
b[13615] == 13615 && 
b[13616] == 13616 && 
b[13617] == 13617 && 
b[13618] == 13618 && 
b[13619] == 13619 && 
b[13620] == 13620 && 
b[13621] == 13621 && 
b[13622] == 13622 && 
b[13623] == 13623 && 
b[13624] == 13624 && 
b[13625] == 13625 && 
b[13626] == 13626 && 
b[13627] == 13627 && 
b[13628] == 13628 && 
b[13629] == 13629 && 
b[13630] == 13630 && 
b[13631] == 13631 && 
b[13632] == 13632 && 
b[13633] == 13633 && 
b[13634] == 13634 && 
b[13635] == 13635 && 
b[13636] == 13636 && 
b[13637] == 13637 && 
b[13638] == 13638 && 
b[13639] == 13639 && 
b[13640] == 13640 && 
b[13641] == 13641 && 
b[13642] == 13642 && 
b[13643] == 13643 && 
b[13644] == 13644 && 
b[13645] == 13645 && 
b[13646] == 13646 && 
b[13647] == 13647 && 
b[13648] == 13648 && 
b[13649] == 13649 && 
b[13650] == 13650 && 
b[13651] == 13651 && 
b[13652] == 13652 && 
b[13653] == 13653 && 
b[13654] == 13654 && 
b[13655] == 13655 && 
b[13656] == 13656 && 
b[13657] == 13657 && 
b[13658] == 13658 && 
b[13659] == 13659 && 
b[13660] == 13660 && 
b[13661] == 13661 && 
b[13662] == 13662 && 
b[13663] == 13663 && 
b[13664] == 13664 && 
b[13665] == 13665 && 
b[13666] == 13666 && 
b[13667] == 13667 && 
b[13668] == 13668 && 
b[13669] == 13669 && 
b[13670] == 13670 && 
b[13671] == 13671 && 
b[13672] == 13672 && 
b[13673] == 13673 && 
b[13674] == 13674 && 
b[13675] == 13675 && 
b[13676] == 13676 && 
b[13677] == 13677 && 
b[13678] == 13678 && 
b[13679] == 13679 && 
b[13680] == 13680 && 
b[13681] == 13681 && 
b[13682] == 13682 && 
b[13683] == 13683 && 
b[13684] == 13684 && 
b[13685] == 13685 && 
b[13686] == 13686 && 
b[13687] == 13687 && 
b[13688] == 13688 && 
b[13689] == 13689 && 
b[13690] == 13690 && 
b[13691] == 13691 && 
b[13692] == 13692 && 
b[13693] == 13693 && 
b[13694] == 13694 && 
b[13695] == 13695 && 
b[13696] == 13696 && 
b[13697] == 13697 && 
b[13698] == 13698 && 
b[13699] == 13699 && 
b[13700] == 13700 && 
b[13701] == 13701 && 
b[13702] == 13702 && 
b[13703] == 13703 && 
b[13704] == 13704 && 
b[13705] == 13705 && 
b[13706] == 13706 && 
b[13707] == 13707 && 
b[13708] == 13708 && 
b[13709] == 13709 && 
b[13710] == 13710 && 
b[13711] == 13711 && 
b[13712] == 13712 && 
b[13713] == 13713 && 
b[13714] == 13714 && 
b[13715] == 13715 && 
b[13716] == 13716 && 
b[13717] == 13717 && 
b[13718] == 13718 && 
b[13719] == 13719 && 
b[13720] == 13720 && 
b[13721] == 13721 && 
b[13722] == 13722 && 
b[13723] == 13723 && 
b[13724] == 13724 && 
b[13725] == 13725 && 
b[13726] == 13726 && 
b[13727] == 13727 && 
b[13728] == 13728 && 
b[13729] == 13729 && 
b[13730] == 13730 && 
b[13731] == 13731 && 
b[13732] == 13732 && 
b[13733] == 13733 && 
b[13734] == 13734 && 
b[13735] == 13735 && 
b[13736] == 13736 && 
b[13737] == 13737 && 
b[13738] == 13738 && 
b[13739] == 13739 && 
b[13740] == 13740 && 
b[13741] == 13741 && 
b[13742] == 13742 && 
b[13743] == 13743 && 
b[13744] == 13744 && 
b[13745] == 13745 && 
b[13746] == 13746 && 
b[13747] == 13747 && 
b[13748] == 13748 && 
b[13749] == 13749 && 
b[13750] == 13750 && 
b[13751] == 13751 && 
b[13752] == 13752 && 
b[13753] == 13753 && 
b[13754] == 13754 && 
b[13755] == 13755 && 
b[13756] == 13756 && 
b[13757] == 13757 && 
b[13758] == 13758 && 
b[13759] == 13759 && 
b[13760] == 13760 && 
b[13761] == 13761 && 
b[13762] == 13762 && 
b[13763] == 13763 && 
b[13764] == 13764 && 
b[13765] == 13765 && 
b[13766] == 13766 && 
b[13767] == 13767 && 
b[13768] == 13768 && 
b[13769] == 13769 && 
b[13770] == 13770 && 
b[13771] == 13771 && 
b[13772] == 13772 && 
b[13773] == 13773 && 
b[13774] == 13774 && 
b[13775] == 13775 && 
b[13776] == 13776 && 
b[13777] == 13777 && 
b[13778] == 13778 && 
b[13779] == 13779 && 
b[13780] == 13780 && 
b[13781] == 13781 && 
b[13782] == 13782 && 
b[13783] == 13783 && 
b[13784] == 13784 && 
b[13785] == 13785 && 
b[13786] == 13786 && 
b[13787] == 13787 && 
b[13788] == 13788 && 
b[13789] == 13789 && 
b[13790] == 13790 && 
b[13791] == 13791 && 
b[13792] == 13792 && 
b[13793] == 13793 && 
b[13794] == 13794 && 
b[13795] == 13795 && 
b[13796] == 13796 && 
b[13797] == 13797 && 
b[13798] == 13798 && 
b[13799] == 13799 && 
b[13800] == 13800 && 
b[13801] == 13801 && 
b[13802] == 13802 && 
b[13803] == 13803 && 
b[13804] == 13804 && 
b[13805] == 13805 && 
b[13806] == 13806 && 
b[13807] == 13807 && 
b[13808] == 13808 && 
b[13809] == 13809 && 
b[13810] == 13810 && 
b[13811] == 13811 && 
b[13812] == 13812 && 
b[13813] == 13813 && 
b[13814] == 13814 && 
b[13815] == 13815 && 
b[13816] == 13816 && 
b[13817] == 13817 && 
b[13818] == 13818 && 
b[13819] == 13819 && 
b[13820] == 13820 && 
b[13821] == 13821 && 
b[13822] == 13822 && 
b[13823] == 13823 && 
b[13824] == 13824 && 
b[13825] == 13825 && 
b[13826] == 13826 && 
b[13827] == 13827 && 
b[13828] == 13828 && 
b[13829] == 13829 && 
b[13830] == 13830 && 
b[13831] == 13831 && 
b[13832] == 13832 && 
b[13833] == 13833 && 
b[13834] == 13834 && 
b[13835] == 13835 && 
b[13836] == 13836 && 
b[13837] == 13837 && 
b[13838] == 13838 && 
b[13839] == 13839 && 
b[13840] == 13840 && 
b[13841] == 13841 && 
b[13842] == 13842 && 
b[13843] == 13843 && 
b[13844] == 13844 && 
b[13845] == 13845 && 
b[13846] == 13846 && 
b[13847] == 13847 && 
b[13848] == 13848 && 
b[13849] == 13849 && 
b[13850] == 13850 && 
b[13851] == 13851 && 
b[13852] == 13852 && 
b[13853] == 13853 && 
b[13854] == 13854 && 
b[13855] == 13855 && 
b[13856] == 13856 && 
b[13857] == 13857 && 
b[13858] == 13858 && 
b[13859] == 13859 && 
b[13860] == 13860 && 
b[13861] == 13861 && 
b[13862] == 13862 && 
b[13863] == 13863 && 
b[13864] == 13864 && 
b[13865] == 13865 && 
b[13866] == 13866 && 
b[13867] == 13867 && 
b[13868] == 13868 && 
b[13869] == 13869 && 
b[13870] == 13870 && 
b[13871] == 13871 && 
b[13872] == 13872 && 
b[13873] == 13873 && 
b[13874] == 13874 && 
b[13875] == 13875 && 
b[13876] == 13876 && 
b[13877] == 13877 && 
b[13878] == 13878 && 
b[13879] == 13879 && 
b[13880] == 13880 && 
b[13881] == 13881 && 
b[13882] == 13882 && 
b[13883] == 13883 && 
b[13884] == 13884 && 
b[13885] == 13885 && 
b[13886] == 13886 && 
b[13887] == 13887 && 
b[13888] == 13888 && 
b[13889] == 13889 && 
b[13890] == 13890 && 
b[13891] == 13891 && 
b[13892] == 13892 && 
b[13893] == 13893 && 
b[13894] == 13894 && 
b[13895] == 13895 && 
b[13896] == 13896 && 
b[13897] == 13897 && 
b[13898] == 13898 && 
b[13899] == 13899 && 
b[13900] == 13900 && 
b[13901] == 13901 && 
b[13902] == 13902 && 
b[13903] == 13903 && 
b[13904] == 13904 && 
b[13905] == 13905 && 
b[13906] == 13906 && 
b[13907] == 13907 && 
b[13908] == 13908 && 
b[13909] == 13909 && 
b[13910] == 13910 && 
b[13911] == 13911 && 
b[13912] == 13912 && 
b[13913] == 13913 && 
b[13914] == 13914 && 
b[13915] == 13915 && 
b[13916] == 13916 && 
b[13917] == 13917 && 
b[13918] == 13918 && 
b[13919] == 13919 && 
b[13920] == 13920 && 
b[13921] == 13921 && 
b[13922] == 13922 && 
b[13923] == 13923 && 
b[13924] == 13924 && 
b[13925] == 13925 && 
b[13926] == 13926 && 
b[13927] == 13927 && 
b[13928] == 13928 && 
b[13929] == 13929 && 
b[13930] == 13930 && 
b[13931] == 13931 && 
b[13932] == 13932 && 
b[13933] == 13933 && 
b[13934] == 13934 && 
b[13935] == 13935 && 
b[13936] == 13936 && 
b[13937] == 13937 && 
b[13938] == 13938 && 
b[13939] == 13939 && 
b[13940] == 13940 && 
b[13941] == 13941 && 
b[13942] == 13942 && 
b[13943] == 13943 && 
b[13944] == 13944 && 
b[13945] == 13945 && 
b[13946] == 13946 && 
b[13947] == 13947 && 
b[13948] == 13948 && 
b[13949] == 13949 && 
b[13950] == 13950 && 
b[13951] == 13951 && 
b[13952] == 13952 && 
b[13953] == 13953 && 
b[13954] == 13954 && 
b[13955] == 13955 && 
b[13956] == 13956 && 
b[13957] == 13957 && 
b[13958] == 13958 && 
b[13959] == 13959 && 
b[13960] == 13960 && 
b[13961] == 13961 && 
b[13962] == 13962 && 
b[13963] == 13963 && 
b[13964] == 13964 && 
b[13965] == 13965 && 
b[13966] == 13966 && 
b[13967] == 13967 && 
b[13968] == 13968 && 
b[13969] == 13969 && 
b[13970] == 13970 && 
b[13971] == 13971 && 
b[13972] == 13972 && 
b[13973] == 13973 && 
b[13974] == 13974 && 
b[13975] == 13975 && 
b[13976] == 13976 && 
b[13977] == 13977 && 
b[13978] == 13978 && 
b[13979] == 13979 && 
b[13980] == 13980 && 
b[13981] == 13981 && 
b[13982] == 13982 && 
b[13983] == 13983 && 
b[13984] == 13984 && 
b[13985] == 13985 && 
b[13986] == 13986 && 
b[13987] == 13987 && 
b[13988] == 13988 && 
b[13989] == 13989 && 
b[13990] == 13990 && 
b[13991] == 13991 && 
b[13992] == 13992 && 
b[13993] == 13993 && 
b[13994] == 13994 && 
b[13995] == 13995 && 
b[13996] == 13996 && 
b[13997] == 13997 && 
b[13998] == 13998 && 
b[13999] == 13999 && 
b[14000] == 14000 && 
b[14001] == 14001 && 
b[14002] == 14002 && 
b[14003] == 14003 && 
b[14004] == 14004 && 
b[14005] == 14005 && 
b[14006] == 14006 && 
b[14007] == 14007 && 
b[14008] == 14008 && 
b[14009] == 14009 && 
b[14010] == 14010 && 
b[14011] == 14011 && 
b[14012] == 14012 && 
b[14013] == 14013 && 
b[14014] == 14014 && 
b[14015] == 14015 && 
b[14016] == 14016 && 
b[14017] == 14017 && 
b[14018] == 14018 && 
b[14019] == 14019 && 
b[14020] == 14020 && 
b[14021] == 14021 && 
b[14022] == 14022 && 
b[14023] == 14023 && 
b[14024] == 14024 && 
b[14025] == 14025 && 
b[14026] == 14026 && 
b[14027] == 14027 && 
b[14028] == 14028 && 
b[14029] == 14029 && 
b[14030] == 14030 && 
b[14031] == 14031 && 
b[14032] == 14032 && 
b[14033] == 14033 && 
b[14034] == 14034 && 
b[14035] == 14035 && 
b[14036] == 14036 && 
b[14037] == 14037 && 
b[14038] == 14038 && 
b[14039] == 14039 && 
b[14040] == 14040 && 
b[14041] == 14041 && 
b[14042] == 14042 && 
b[14043] == 14043 && 
b[14044] == 14044 && 
b[14045] == 14045 && 
b[14046] == 14046 && 
b[14047] == 14047 && 
b[14048] == 14048 && 
b[14049] == 14049 && 
b[14050] == 14050 && 
b[14051] == 14051 && 
b[14052] == 14052 && 
b[14053] == 14053 && 
b[14054] == 14054 && 
b[14055] == 14055 && 
b[14056] == 14056 && 
b[14057] == 14057 && 
b[14058] == 14058 && 
b[14059] == 14059 && 
b[14060] == 14060 && 
b[14061] == 14061 && 
b[14062] == 14062 && 
b[14063] == 14063 && 
b[14064] == 14064 && 
b[14065] == 14065 && 
b[14066] == 14066 && 
b[14067] == 14067 && 
b[14068] == 14068 && 
b[14069] == 14069 && 
b[14070] == 14070 && 
b[14071] == 14071 && 
b[14072] == 14072 && 
b[14073] == 14073 && 
b[14074] == 14074 && 
b[14075] == 14075 && 
b[14076] == 14076 && 
b[14077] == 14077 && 
b[14078] == 14078 && 
b[14079] == 14079 && 
b[14080] == 14080 && 
b[14081] == 14081 && 
b[14082] == 14082 && 
b[14083] == 14083 && 
b[14084] == 14084 && 
b[14085] == 14085 && 
b[14086] == 14086 && 
b[14087] == 14087 && 
b[14088] == 14088 && 
b[14089] == 14089 && 
b[14090] == 14090 && 
b[14091] == 14091 && 
b[14092] == 14092 && 
b[14093] == 14093 && 
b[14094] == 14094 && 
b[14095] == 14095 && 
b[14096] == 14096 && 
b[14097] == 14097 && 
b[14098] == 14098 && 
b[14099] == 14099 && 
b[14100] == 14100 && 
b[14101] == 14101 && 
b[14102] == 14102 && 
b[14103] == 14103 && 
b[14104] == 14104 && 
b[14105] == 14105 && 
b[14106] == 14106 && 
b[14107] == 14107 && 
b[14108] == 14108 && 
b[14109] == 14109 && 
b[14110] == 14110 && 
b[14111] == 14111 && 
b[14112] == 14112 && 
b[14113] == 14113 && 
b[14114] == 14114 && 
b[14115] == 14115 && 
b[14116] == 14116 && 
b[14117] == 14117 && 
b[14118] == 14118 && 
b[14119] == 14119 && 
b[14120] == 14120 && 
b[14121] == 14121 && 
b[14122] == 14122 && 
b[14123] == 14123 && 
b[14124] == 14124 && 
b[14125] == 14125 && 
b[14126] == 14126 && 
b[14127] == 14127 && 
b[14128] == 14128 && 
b[14129] == 14129 && 
b[14130] == 14130 && 
b[14131] == 14131 && 
b[14132] == 14132 && 
b[14133] == 14133 && 
b[14134] == 14134 && 
b[14135] == 14135 && 
b[14136] == 14136 && 
b[14137] == 14137 && 
b[14138] == 14138 && 
b[14139] == 14139 && 
b[14140] == 14140 && 
b[14141] == 14141 && 
b[14142] == 14142 && 
b[14143] == 14143 && 
b[14144] == 14144 && 
b[14145] == 14145 && 
b[14146] == 14146 && 
b[14147] == 14147 && 
b[14148] == 14148 && 
b[14149] == 14149 && 
b[14150] == 14150 && 
b[14151] == 14151 && 
b[14152] == 14152 && 
b[14153] == 14153 && 
b[14154] == 14154 && 
b[14155] == 14155 && 
b[14156] == 14156 && 
b[14157] == 14157 && 
b[14158] == 14158 && 
b[14159] == 14159 && 
b[14160] == 14160 && 
b[14161] == 14161 && 
b[14162] == 14162 && 
b[14163] == 14163 && 
b[14164] == 14164 && 
b[14165] == 14165 && 
b[14166] == 14166 && 
b[14167] == 14167 && 
b[14168] == 14168 && 
b[14169] == 14169 && 
b[14170] == 14170 && 
b[14171] == 14171 && 
b[14172] == 14172 && 
b[14173] == 14173 && 
b[14174] == 14174 && 
b[14175] == 14175 && 
b[14176] == 14176 && 
b[14177] == 14177 && 
b[14178] == 14178 && 
b[14179] == 14179 && 
b[14180] == 14180 && 
b[14181] == 14181 && 
b[14182] == 14182 && 
b[14183] == 14183 && 
b[14184] == 14184 && 
b[14185] == 14185 && 
b[14186] == 14186 && 
b[14187] == 14187 && 
b[14188] == 14188 && 
b[14189] == 14189 && 
b[14190] == 14190 && 
b[14191] == 14191 && 
b[14192] == 14192 && 
b[14193] == 14193 && 
b[14194] == 14194 && 
b[14195] == 14195 && 
b[14196] == 14196 && 
b[14197] == 14197 && 
b[14198] == 14198 && 
b[14199] == 14199 && 
b[14200] == 14200 && 
b[14201] == 14201 && 
b[14202] == 14202 && 
b[14203] == 14203 && 
b[14204] == 14204 && 
b[14205] == 14205 && 
b[14206] == 14206 && 
b[14207] == 14207 && 
b[14208] == 14208 && 
b[14209] == 14209 && 
b[14210] == 14210 && 
b[14211] == 14211 && 
b[14212] == 14212 && 
b[14213] == 14213 && 
b[14214] == 14214 && 
b[14215] == 14215 && 
b[14216] == 14216 && 
b[14217] == 14217 && 
b[14218] == 14218 && 
b[14219] == 14219 && 
b[14220] == 14220 && 
b[14221] == 14221 && 
b[14222] == 14222 && 
b[14223] == 14223 && 
b[14224] == 14224 && 
b[14225] == 14225 && 
b[14226] == 14226 && 
b[14227] == 14227 && 
b[14228] == 14228 && 
b[14229] == 14229 && 
b[14230] == 14230 && 
b[14231] == 14231 && 
b[14232] == 14232 && 
b[14233] == 14233 && 
b[14234] == 14234 && 
b[14235] == 14235 && 
b[14236] == 14236 && 
b[14237] == 14237 && 
b[14238] == 14238 && 
b[14239] == 14239 && 
b[14240] == 14240 && 
b[14241] == 14241 && 
b[14242] == 14242 && 
b[14243] == 14243 && 
b[14244] == 14244 && 
b[14245] == 14245 && 
b[14246] == 14246 && 
b[14247] == 14247 && 
b[14248] == 14248 && 
b[14249] == 14249 && 
b[14250] == 14250 && 
b[14251] == 14251 && 
b[14252] == 14252 && 
b[14253] == 14253 && 
b[14254] == 14254 && 
b[14255] == 14255 && 
b[14256] == 14256 && 
b[14257] == 14257 && 
b[14258] == 14258 && 
b[14259] == 14259 && 
b[14260] == 14260 && 
b[14261] == 14261 && 
b[14262] == 14262 && 
b[14263] == 14263 && 
b[14264] == 14264 && 
b[14265] == 14265 && 
b[14266] == 14266 && 
b[14267] == 14267 && 
b[14268] == 14268 && 
b[14269] == 14269 && 
b[14270] == 14270 && 
b[14271] == 14271 && 
b[14272] == 14272 && 
b[14273] == 14273 && 
b[14274] == 14274 && 
b[14275] == 14275 && 
b[14276] == 14276 && 
b[14277] == 14277 && 
b[14278] == 14278 && 
b[14279] == 14279 && 
b[14280] == 14280 && 
b[14281] == 14281 && 
b[14282] == 14282 && 
b[14283] == 14283 && 
b[14284] == 14284 && 
b[14285] == 14285 && 
b[14286] == 14286 && 
b[14287] == 14287 && 
b[14288] == 14288 && 
b[14289] == 14289 && 
b[14290] == 14290 && 
b[14291] == 14291 && 
b[14292] == 14292 && 
b[14293] == 14293 && 
b[14294] == 14294 && 
b[14295] == 14295 && 
b[14296] == 14296 && 
b[14297] == 14297 && 
b[14298] == 14298 && 
b[14299] == 14299 && 
b[14300] == 14300 && 
b[14301] == 14301 && 
b[14302] == 14302 && 
b[14303] == 14303 && 
b[14304] == 14304 && 
b[14305] == 14305 && 
b[14306] == 14306 && 
b[14307] == 14307 && 
b[14308] == 14308 && 
b[14309] == 14309 && 
b[14310] == 14310 && 
b[14311] == 14311 && 
b[14312] == 14312 && 
b[14313] == 14313 && 
b[14314] == 14314 && 
b[14315] == 14315 && 
b[14316] == 14316 && 
b[14317] == 14317 && 
b[14318] == 14318 && 
b[14319] == 14319 && 
b[14320] == 14320 && 
b[14321] == 14321 && 
b[14322] == 14322 && 
b[14323] == 14323 && 
b[14324] == 14324 && 
b[14325] == 14325 && 
b[14326] == 14326 && 
b[14327] == 14327 && 
b[14328] == 14328 && 
b[14329] == 14329 && 
b[14330] == 14330 && 
b[14331] == 14331 && 
b[14332] == 14332 && 
b[14333] == 14333 && 
b[14334] == 14334 && 
b[14335] == 14335 && 
b[14336] == 14336 && 
b[14337] == 14337 && 
b[14338] == 14338 && 
b[14339] == 14339 && 
b[14340] == 14340 && 
b[14341] == 14341 && 
b[14342] == 14342 && 
b[14343] == 14343 && 
b[14344] == 14344 && 
b[14345] == 14345 && 
b[14346] == 14346 && 
b[14347] == 14347 && 
b[14348] == 14348 && 
b[14349] == 14349 && 
b[14350] == 14350 && 
b[14351] == 14351 && 
b[14352] == 14352 && 
b[14353] == 14353 && 
b[14354] == 14354 && 
b[14355] == 14355 && 
b[14356] == 14356 && 
b[14357] == 14357 && 
b[14358] == 14358 && 
b[14359] == 14359 && 
b[14360] == 14360 && 
b[14361] == 14361 && 
b[14362] == 14362 && 
b[14363] == 14363 && 
b[14364] == 14364 && 
b[14365] == 14365 && 
b[14366] == 14366 && 
b[14367] == 14367 && 
b[14368] == 14368 && 
b[14369] == 14369 && 
b[14370] == 14370 && 
b[14371] == 14371 && 
b[14372] == 14372 && 
b[14373] == 14373 && 
b[14374] == 14374 && 
b[14375] == 14375 && 
b[14376] == 14376 && 
b[14377] == 14377 && 
b[14378] == 14378 && 
b[14379] == 14379 && 
b[14380] == 14380 && 
b[14381] == 14381 && 
b[14382] == 14382 && 
b[14383] == 14383 && 
b[14384] == 14384 && 
b[14385] == 14385 && 
b[14386] == 14386 && 
b[14387] == 14387 && 
b[14388] == 14388 && 
b[14389] == 14389 && 
b[14390] == 14390 && 
b[14391] == 14391 && 
b[14392] == 14392 && 
b[14393] == 14393 && 
b[14394] == 14394 && 
b[14395] == 14395 && 
b[14396] == 14396 && 
b[14397] == 14397 && 
b[14398] == 14398 && 
b[14399] == 14399 && 
b[14400] == 14400 && 
b[14401] == 14401 && 
b[14402] == 14402 && 
b[14403] == 14403 && 
b[14404] == 14404 && 
b[14405] == 14405 && 
b[14406] == 14406 && 
b[14407] == 14407 && 
b[14408] == 14408 && 
b[14409] == 14409 && 
b[14410] == 14410 && 
b[14411] == 14411 && 
b[14412] == 14412 && 
b[14413] == 14413 && 
b[14414] == 14414 && 
b[14415] == 14415 && 
b[14416] == 14416 && 
b[14417] == 14417 && 
b[14418] == 14418 && 
b[14419] == 14419 && 
b[14420] == 14420 && 
b[14421] == 14421 && 
b[14422] == 14422 && 
b[14423] == 14423 && 
b[14424] == 14424 && 
b[14425] == 14425 && 
b[14426] == 14426 && 
b[14427] == 14427 && 
b[14428] == 14428 && 
b[14429] == 14429 && 
b[14430] == 14430 && 
b[14431] == 14431 && 
b[14432] == 14432 && 
b[14433] == 14433 && 
b[14434] == 14434 && 
b[14435] == 14435 && 
b[14436] == 14436 && 
b[14437] == 14437 && 
b[14438] == 14438 && 
b[14439] == 14439 && 
b[14440] == 14440 && 
b[14441] == 14441 && 
b[14442] == 14442 && 
b[14443] == 14443 && 
b[14444] == 14444 && 
b[14445] == 14445 && 
b[14446] == 14446 && 
b[14447] == 14447 && 
b[14448] == 14448 && 
b[14449] == 14449 && 
b[14450] == 14450 && 
b[14451] == 14451 && 
b[14452] == 14452 && 
b[14453] == 14453 && 
b[14454] == 14454 && 
b[14455] == 14455 && 
b[14456] == 14456 && 
b[14457] == 14457 && 
b[14458] == 14458 && 
b[14459] == 14459 && 
b[14460] == 14460 && 
b[14461] == 14461 && 
b[14462] == 14462 && 
b[14463] == 14463 && 
b[14464] == 14464 && 
b[14465] == 14465 && 
b[14466] == 14466 && 
b[14467] == 14467 && 
b[14468] == 14468 && 
b[14469] == 14469 && 
b[14470] == 14470 && 
b[14471] == 14471 && 
b[14472] == 14472 && 
b[14473] == 14473 && 
b[14474] == 14474 && 
b[14475] == 14475 && 
b[14476] == 14476 && 
b[14477] == 14477 && 
b[14478] == 14478 && 
b[14479] == 14479 && 
b[14480] == 14480 && 
b[14481] == 14481 && 
b[14482] == 14482 && 
b[14483] == 14483 && 
b[14484] == 14484 && 
b[14485] == 14485 && 
b[14486] == 14486 && 
b[14487] == 14487 && 
b[14488] == 14488 && 
b[14489] == 14489 && 
b[14490] == 14490 && 
b[14491] == 14491 && 
b[14492] == 14492 && 
b[14493] == 14493 && 
b[14494] == 14494 && 
b[14495] == 14495 && 
b[14496] == 14496 && 
b[14497] == 14497 && 
b[14498] == 14498 && 
b[14499] == 14499 && 
b[14500] == 14500 && 
b[14501] == 14501 && 
b[14502] == 14502 && 
b[14503] == 14503 && 
b[14504] == 14504 && 
b[14505] == 14505 && 
b[14506] == 14506 && 
b[14507] == 14507 && 
b[14508] == 14508 && 
b[14509] == 14509 && 
b[14510] == 14510 && 
b[14511] == 14511 && 
b[14512] == 14512 && 
b[14513] == 14513 && 
b[14514] == 14514 && 
b[14515] == 14515 && 
b[14516] == 14516 && 
b[14517] == 14517 && 
b[14518] == 14518 && 
b[14519] == 14519 && 
b[14520] == 14520 && 
b[14521] == 14521 && 
b[14522] == 14522 && 
b[14523] == 14523 && 
b[14524] == 14524 && 
b[14525] == 14525 && 
b[14526] == 14526 && 
b[14527] == 14527 && 
b[14528] == 14528 && 
b[14529] == 14529 && 
b[14530] == 14530 && 
b[14531] == 14531 && 
b[14532] == 14532 && 
b[14533] == 14533 && 
b[14534] == 14534 && 
b[14535] == 14535 && 
b[14536] == 14536 && 
b[14537] == 14537 && 
b[14538] == 14538 && 
b[14539] == 14539 && 
b[14540] == 14540 && 
b[14541] == 14541 && 
b[14542] == 14542 && 
b[14543] == 14543 && 
b[14544] == 14544 && 
b[14545] == 14545 && 
b[14546] == 14546 && 
b[14547] == 14547 && 
b[14548] == 14548 && 
b[14549] == 14549 && 
b[14550] == 14550 && 
b[14551] == 14551 && 
b[14552] == 14552 && 
b[14553] == 14553 && 
b[14554] == 14554 && 
b[14555] == 14555 && 
b[14556] == 14556 && 
b[14557] == 14557 && 
b[14558] == 14558 && 
b[14559] == 14559 && 
b[14560] == 14560 && 
b[14561] == 14561 && 
b[14562] == 14562 && 
b[14563] == 14563 && 
b[14564] == 14564 && 
b[14565] == 14565 && 
b[14566] == 14566 && 
b[14567] == 14567 && 
b[14568] == 14568 && 
b[14569] == 14569 && 
b[14570] == 14570 && 
b[14571] == 14571 && 
b[14572] == 14572 && 
b[14573] == 14573 && 
b[14574] == 14574 && 
b[14575] == 14575 && 
b[14576] == 14576 && 
b[14577] == 14577 && 
b[14578] == 14578 && 
b[14579] == 14579 && 
b[14580] == 14580 && 
b[14581] == 14581 && 
b[14582] == 14582 && 
b[14583] == 14583 && 
b[14584] == 14584 && 
b[14585] == 14585 && 
b[14586] == 14586 && 
b[14587] == 14587 && 
b[14588] == 14588 && 
b[14589] == 14589 && 
b[14590] == 14590 && 
b[14591] == 14591 && 
b[14592] == 14592 && 
b[14593] == 14593 && 
b[14594] == 14594 && 
b[14595] == 14595 && 
b[14596] == 14596 && 
b[14597] == 14597 && 
b[14598] == 14598 && 
b[14599] == 14599 && 
b[14600] == 14600 && 
b[14601] == 14601 && 
b[14602] == 14602 && 
b[14603] == 14603 && 
b[14604] == 14604 && 
b[14605] == 14605 && 
b[14606] == 14606 && 
b[14607] == 14607 && 
b[14608] == 14608 && 
b[14609] == 14609 && 
b[14610] == 14610 && 
b[14611] == 14611 && 
b[14612] == 14612 && 
b[14613] == 14613 && 
b[14614] == 14614 && 
b[14615] == 14615 && 
b[14616] == 14616 && 
b[14617] == 14617 && 
b[14618] == 14618 && 
b[14619] == 14619 && 
b[14620] == 14620 && 
b[14621] == 14621 && 
b[14622] == 14622 && 
b[14623] == 14623 && 
b[14624] == 14624 && 
b[14625] == 14625 && 
b[14626] == 14626 && 
b[14627] == 14627 && 
b[14628] == 14628 && 
b[14629] == 14629 && 
b[14630] == 14630 && 
b[14631] == 14631 && 
b[14632] == 14632 && 
b[14633] == 14633 && 
b[14634] == 14634 && 
b[14635] == 14635 && 
b[14636] == 14636 && 
b[14637] == 14637 && 
b[14638] == 14638 && 
b[14639] == 14639 && 
b[14640] == 14640 && 
b[14641] == 14641 && 
b[14642] == 14642 && 
b[14643] == 14643 && 
b[14644] == 14644 && 
b[14645] == 14645 && 
b[14646] == 14646 && 
b[14647] == 14647 && 
b[14648] == 14648 && 
b[14649] == 14649 && 
b[14650] == 14650 && 
b[14651] == 14651 && 
b[14652] == 14652 && 
b[14653] == 14653 && 
b[14654] == 14654 && 
b[14655] == 14655 && 
b[14656] == 14656 && 
b[14657] == 14657 && 
b[14658] == 14658 && 
b[14659] == 14659 && 
b[14660] == 14660 && 
b[14661] == 14661 && 
b[14662] == 14662 && 
b[14663] == 14663 && 
b[14664] == 14664 && 
b[14665] == 14665 && 
b[14666] == 14666 && 
b[14667] == 14667 && 
b[14668] == 14668 && 
b[14669] == 14669 && 
b[14670] == 14670 && 
b[14671] == 14671 && 
b[14672] == 14672 && 
b[14673] == 14673 && 
b[14674] == 14674 && 
b[14675] == 14675 && 
b[14676] == 14676 && 
b[14677] == 14677 && 
b[14678] == 14678 && 
b[14679] == 14679 && 
b[14680] == 14680 && 
b[14681] == 14681 && 
b[14682] == 14682 && 
b[14683] == 14683 && 
b[14684] == 14684 && 
b[14685] == 14685 && 
b[14686] == 14686 && 
b[14687] == 14687 && 
b[14688] == 14688 && 
b[14689] == 14689 && 
b[14690] == 14690 && 
b[14691] == 14691 && 
b[14692] == 14692 && 
b[14693] == 14693 && 
b[14694] == 14694 && 
b[14695] == 14695 && 
b[14696] == 14696 && 
b[14697] == 14697 && 
b[14698] == 14698 && 
b[14699] == 14699 && 
b[14700] == 14700 && 
b[14701] == 14701 && 
b[14702] == 14702 && 
b[14703] == 14703 && 
b[14704] == 14704 && 
b[14705] == 14705 && 
b[14706] == 14706 && 
b[14707] == 14707 && 
b[14708] == 14708 && 
b[14709] == 14709 && 
b[14710] == 14710 && 
b[14711] == 14711 && 
b[14712] == 14712 && 
b[14713] == 14713 && 
b[14714] == 14714 && 
b[14715] == 14715 && 
b[14716] == 14716 && 
b[14717] == 14717 && 
b[14718] == 14718 && 
b[14719] == 14719 && 
b[14720] == 14720 && 
b[14721] == 14721 && 
b[14722] == 14722 && 
b[14723] == 14723 && 
b[14724] == 14724 && 
b[14725] == 14725 && 
b[14726] == 14726 && 
b[14727] == 14727 && 
b[14728] == 14728 && 
b[14729] == 14729 && 
b[14730] == 14730 && 
b[14731] == 14731 && 
b[14732] == 14732 && 
b[14733] == 14733 && 
b[14734] == 14734 && 
b[14735] == 14735 && 
b[14736] == 14736 && 
b[14737] == 14737 && 
b[14738] == 14738 && 
b[14739] == 14739 && 
b[14740] == 14740 && 
b[14741] == 14741 && 
b[14742] == 14742 && 
b[14743] == 14743 && 
b[14744] == 14744 && 
b[14745] == 14745 && 
b[14746] == 14746 && 
b[14747] == 14747 && 
b[14748] == 14748 && 
b[14749] == 14749 && 
b[14750] == 14750 && 
b[14751] == 14751 && 
b[14752] == 14752 && 
b[14753] == 14753 && 
b[14754] == 14754 && 
b[14755] == 14755 && 
b[14756] == 14756 && 
b[14757] == 14757 && 
b[14758] == 14758 && 
b[14759] == 14759 && 
b[14760] == 14760 && 
b[14761] == 14761 && 
b[14762] == 14762 && 
b[14763] == 14763 && 
b[14764] == 14764 && 
b[14765] == 14765 && 
b[14766] == 14766 && 
b[14767] == 14767 && 
b[14768] == 14768 && 
b[14769] == 14769 && 
b[14770] == 14770 && 
b[14771] == 14771 && 
b[14772] == 14772 && 
b[14773] == 14773 && 
b[14774] == 14774 && 
b[14775] == 14775 && 
b[14776] == 14776 && 
b[14777] == 14777 && 
b[14778] == 14778 && 
b[14779] == 14779 && 
b[14780] == 14780 && 
b[14781] == 14781 && 
b[14782] == 14782 && 
b[14783] == 14783 && 
b[14784] == 14784 && 
b[14785] == 14785 && 
b[14786] == 14786 && 
b[14787] == 14787 && 
b[14788] == 14788 && 
b[14789] == 14789 && 
b[14790] == 14790 && 
b[14791] == 14791 && 
b[14792] == 14792 && 
b[14793] == 14793 && 
b[14794] == 14794 && 
b[14795] == 14795 && 
b[14796] == 14796 && 
b[14797] == 14797 && 
b[14798] == 14798 && 
b[14799] == 14799 && 
b[14800] == 14800 && 
b[14801] == 14801 && 
b[14802] == 14802 && 
b[14803] == 14803 && 
b[14804] == 14804 && 
b[14805] == 14805 && 
b[14806] == 14806 && 
b[14807] == 14807 && 
b[14808] == 14808 && 
b[14809] == 14809 && 
b[14810] == 14810 && 
b[14811] == 14811 && 
b[14812] == 14812 && 
b[14813] == 14813 && 
b[14814] == 14814 && 
b[14815] == 14815 && 
b[14816] == 14816 && 
b[14817] == 14817 && 
b[14818] == 14818 && 
b[14819] == 14819 && 
b[14820] == 14820 && 
b[14821] == 14821 && 
b[14822] == 14822 && 
b[14823] == 14823 && 
b[14824] == 14824 && 
b[14825] == 14825 && 
b[14826] == 14826 && 
b[14827] == 14827 && 
b[14828] == 14828 && 
b[14829] == 14829 && 
b[14830] == 14830 && 
b[14831] == 14831 && 
b[14832] == 14832 && 
b[14833] == 14833 && 
b[14834] == 14834 && 
b[14835] == 14835 && 
b[14836] == 14836 && 
b[14837] == 14837 && 
b[14838] == 14838 && 
b[14839] == 14839 && 
b[14840] == 14840 && 
b[14841] == 14841 && 
b[14842] == 14842 && 
b[14843] == 14843 && 
b[14844] == 14844 && 
b[14845] == 14845 && 
b[14846] == 14846 && 
b[14847] == 14847 && 
b[14848] == 14848 && 
b[14849] == 14849 && 
b[14850] == 14850 && 
b[14851] == 14851 && 
b[14852] == 14852 && 
b[14853] == 14853 && 
b[14854] == 14854 && 
b[14855] == 14855 && 
b[14856] == 14856 && 
b[14857] == 14857 && 
b[14858] == 14858 && 
b[14859] == 14859 && 
b[14860] == 14860 && 
b[14861] == 14861 && 
b[14862] == 14862 && 
b[14863] == 14863 && 
b[14864] == 14864 && 
b[14865] == 14865 && 
b[14866] == 14866 && 
b[14867] == 14867 && 
b[14868] == 14868 && 
b[14869] == 14869 && 
b[14870] == 14870 && 
b[14871] == 14871 && 
b[14872] == 14872 && 
b[14873] == 14873 && 
b[14874] == 14874 && 
b[14875] == 14875 && 
b[14876] == 14876 && 
b[14877] == 14877 && 
b[14878] == 14878 && 
b[14879] == 14879 && 
b[14880] == 14880 && 
b[14881] == 14881 && 
b[14882] == 14882 && 
b[14883] == 14883 && 
b[14884] == 14884 && 
b[14885] == 14885 && 
b[14886] == 14886 && 
b[14887] == 14887 && 
b[14888] == 14888 && 
b[14889] == 14889 && 
b[14890] == 14890 && 
b[14891] == 14891 && 
b[14892] == 14892 && 
b[14893] == 14893 && 
b[14894] == 14894 && 
b[14895] == 14895 && 
b[14896] == 14896 && 
b[14897] == 14897 && 
b[14898] == 14898 && 
b[14899] == 14899 && 
b[14900] == 14900 && 
b[14901] == 14901 && 
b[14902] == 14902 && 
b[14903] == 14903 && 
b[14904] == 14904 && 
b[14905] == 14905 && 
b[14906] == 14906 && 
b[14907] == 14907 && 
b[14908] == 14908 && 
b[14909] == 14909 && 
b[14910] == 14910 && 
b[14911] == 14911 && 
b[14912] == 14912 && 
b[14913] == 14913 && 
b[14914] == 14914 && 
b[14915] == 14915 && 
b[14916] == 14916 && 
b[14917] == 14917 && 
b[14918] == 14918 && 
b[14919] == 14919 && 
b[14920] == 14920 && 
b[14921] == 14921 && 
b[14922] == 14922 && 
b[14923] == 14923 && 
b[14924] == 14924 && 
b[14925] == 14925 && 
b[14926] == 14926 && 
b[14927] == 14927 && 
b[14928] == 14928 && 
b[14929] == 14929 && 
b[14930] == 14930 && 
b[14931] == 14931 && 
b[14932] == 14932 && 
b[14933] == 14933 && 
b[14934] == 14934 && 
b[14935] == 14935 && 
b[14936] == 14936 && 
b[14937] == 14937 && 
b[14938] == 14938 && 
b[14939] == 14939 && 
b[14940] == 14940 && 
b[14941] == 14941 && 
b[14942] == 14942 && 
b[14943] == 14943 && 
b[14944] == 14944 && 
b[14945] == 14945 && 
b[14946] == 14946 && 
b[14947] == 14947 && 
b[14948] == 14948 && 
b[14949] == 14949 && 
b[14950] == 14950 && 
b[14951] == 14951 && 
b[14952] == 14952 && 
b[14953] == 14953 && 
b[14954] == 14954 && 
b[14955] == 14955 && 
b[14956] == 14956 && 
b[14957] == 14957 && 
b[14958] == 14958 && 
b[14959] == 14959 && 
b[14960] == 14960 && 
b[14961] == 14961 && 
b[14962] == 14962 && 
b[14963] == 14963 && 
b[14964] == 14964 && 
b[14965] == 14965 && 
b[14966] == 14966 && 
b[14967] == 14967 && 
b[14968] == 14968 && 
b[14969] == 14969 && 
b[14970] == 14970 && 
b[14971] == 14971 && 
b[14972] == 14972 && 
b[14973] == 14973 && 
b[14974] == 14974 && 
b[14975] == 14975 && 
b[14976] == 14976 && 
b[14977] == 14977 && 
b[14978] == 14978 && 
b[14979] == 14979 && 
b[14980] == 14980 && 
b[14981] == 14981 && 
b[14982] == 14982 && 
b[14983] == 14983 && 
b[14984] == 14984 && 
b[14985] == 14985 && 
b[14986] == 14986 && 
b[14987] == 14987 && 
b[14988] == 14988 && 
b[14989] == 14989 && 
b[14990] == 14990 && 
b[14991] == 14991 && 
b[14992] == 14992 && 
b[14993] == 14993 && 
b[14994] == 14994 && 
b[14995] == 14995 && 
b[14996] == 14996 && 
b[14997] == 14997 && 
b[14998] == 14998 && 
b[14999] == 14999 && 
b[15000] == 15000 && 
b[15001] == 15001 && 
b[15002] == 15002 && 
b[15003] == 15003 && 
b[15004] == 15004 && 
b[15005] == 15005 && 
b[15006] == 15006 && 
b[15007] == 15007 && 
b[15008] == 15008 && 
b[15009] == 15009 && 
b[15010] == 15010 && 
b[15011] == 15011 && 
b[15012] == 15012 && 
b[15013] == 15013 && 
b[15014] == 15014 && 
b[15015] == 15015 && 
b[15016] == 15016 && 
b[15017] == 15017 && 
b[15018] == 15018 && 
b[15019] == 15019 && 
b[15020] == 15020 && 
b[15021] == 15021 && 
b[15022] == 15022 && 
b[15023] == 15023 && 
b[15024] == 15024 && 
b[15025] == 15025 && 
b[15026] == 15026 && 
b[15027] == 15027 && 
b[15028] == 15028 && 
b[15029] == 15029 && 
b[15030] == 15030 && 
b[15031] == 15031 && 
b[15032] == 15032 && 
b[15033] == 15033 && 
b[15034] == 15034 && 
b[15035] == 15035 && 
b[15036] == 15036 && 
b[15037] == 15037 && 
b[15038] == 15038 && 
b[15039] == 15039 && 
b[15040] == 15040 && 
b[15041] == 15041 && 
b[15042] == 15042 && 
b[15043] == 15043 && 
b[15044] == 15044 && 
b[15045] == 15045 && 
b[15046] == 15046 && 
b[15047] == 15047 && 
b[15048] == 15048 && 
b[15049] == 15049 && 
b[15050] == 15050 && 
b[15051] == 15051 && 
b[15052] == 15052 && 
b[15053] == 15053 && 
b[15054] == 15054 && 
b[15055] == 15055 && 
b[15056] == 15056 && 
b[15057] == 15057 && 
b[15058] == 15058 && 
b[15059] == 15059 && 
b[15060] == 15060 && 
b[15061] == 15061 && 
b[15062] == 15062 && 
b[15063] == 15063 && 
b[15064] == 15064 && 
b[15065] == 15065 && 
b[15066] == 15066 && 
b[15067] == 15067 && 
b[15068] == 15068 && 
b[15069] == 15069 && 
b[15070] == 15070 && 
b[15071] == 15071 && 
b[15072] == 15072 && 
b[15073] == 15073 && 
b[15074] == 15074 && 
b[15075] == 15075 && 
b[15076] == 15076 && 
b[15077] == 15077 && 
b[15078] == 15078 && 
b[15079] == 15079 && 
b[15080] == 15080 && 
b[15081] == 15081 && 
b[15082] == 15082 && 
b[15083] == 15083 && 
b[15084] == 15084 && 
b[15085] == 15085 && 
b[15086] == 15086 && 
b[15087] == 15087 && 
b[15088] == 15088 && 
b[15089] == 15089 && 
b[15090] == 15090 && 
b[15091] == 15091 && 
b[15092] == 15092 && 
b[15093] == 15093 && 
b[15094] == 15094 && 
b[15095] == 15095 && 
b[15096] == 15096 && 
b[15097] == 15097 && 
b[15098] == 15098 && 
b[15099] == 15099 && 
b[15100] == 15100 && 
b[15101] == 15101 && 
b[15102] == 15102 && 
b[15103] == 15103 && 
b[15104] == 15104 && 
b[15105] == 15105 && 
b[15106] == 15106 && 
b[15107] == 15107 && 
b[15108] == 15108 && 
b[15109] == 15109 && 
b[15110] == 15110 && 
b[15111] == 15111 && 
b[15112] == 15112 && 
b[15113] == 15113 && 
b[15114] == 15114 && 
b[15115] == 15115 && 
b[15116] == 15116 && 
b[15117] == 15117 && 
b[15118] == 15118 && 
b[15119] == 15119 && 
b[15120] == 15120 && 
b[15121] == 15121 && 
b[15122] == 15122 && 
b[15123] == 15123 && 
b[15124] == 15124 && 
b[15125] == 15125 && 
b[15126] == 15126 && 
b[15127] == 15127 && 
b[15128] == 15128 && 
b[15129] == 15129 && 
b[15130] == 15130 && 
b[15131] == 15131 && 
b[15132] == 15132 && 
b[15133] == 15133 && 
b[15134] == 15134 && 
b[15135] == 15135 && 
b[15136] == 15136 && 
b[15137] == 15137 && 
b[15138] == 15138 && 
b[15139] == 15139 && 
b[15140] == 15140 && 
b[15141] == 15141 && 
b[15142] == 15142 && 
b[15143] == 15143 && 
b[15144] == 15144 && 
b[15145] == 15145 && 
b[15146] == 15146 && 
b[15147] == 15147 && 
b[15148] == 15148 && 
b[15149] == 15149 && 
b[15150] == 15150 && 
b[15151] == 15151 && 
b[15152] == 15152 && 
b[15153] == 15153 && 
b[15154] == 15154 && 
b[15155] == 15155 && 
b[15156] == 15156 && 
b[15157] == 15157 && 
b[15158] == 15158 && 
b[15159] == 15159 && 
b[15160] == 15160 && 
b[15161] == 15161 && 
b[15162] == 15162 && 
b[15163] == 15163 && 
b[15164] == 15164 && 
b[15165] == 15165 && 
b[15166] == 15166 && 
b[15167] == 15167 && 
b[15168] == 15168 && 
b[15169] == 15169 && 
b[15170] == 15170 && 
b[15171] == 15171 && 
b[15172] == 15172 && 
b[15173] == 15173 && 
b[15174] == 15174 && 
b[15175] == 15175 && 
b[15176] == 15176 && 
b[15177] == 15177 && 
b[15178] == 15178 && 
b[15179] == 15179 && 
b[15180] == 15180 && 
b[15181] == 15181 && 
b[15182] == 15182 && 
b[15183] == 15183 && 
b[15184] == 15184 && 
b[15185] == 15185 && 
b[15186] == 15186 && 
b[15187] == 15187 && 
b[15188] == 15188 && 
b[15189] == 15189 && 
b[15190] == 15190 && 
b[15191] == 15191 && 
b[15192] == 15192 && 
b[15193] == 15193 && 
b[15194] == 15194 && 
b[15195] == 15195 && 
b[15196] == 15196 && 
b[15197] == 15197 && 
b[15198] == 15198 && 
b[15199] == 15199 && 
b[15200] == 15200 && 
b[15201] == 15201 && 
b[15202] == 15202 && 
b[15203] == 15203 && 
b[15204] == 15204 && 
b[15205] == 15205 && 
b[15206] == 15206 && 
b[15207] == 15207 && 
b[15208] == 15208 && 
b[15209] == 15209 && 
b[15210] == 15210 && 
b[15211] == 15211 && 
b[15212] == 15212 && 
b[15213] == 15213 && 
b[15214] == 15214 && 
b[15215] == 15215 && 
b[15216] == 15216 && 
b[15217] == 15217 && 
b[15218] == 15218 && 
b[15219] == 15219 && 
b[15220] == 15220 && 
b[15221] == 15221 && 
b[15222] == 15222 && 
b[15223] == 15223 && 
b[15224] == 15224 && 
b[15225] == 15225 && 
b[15226] == 15226 && 
b[15227] == 15227 && 
b[15228] == 15228 && 
b[15229] == 15229 && 
b[15230] == 15230 && 
b[15231] == 15231 && 
b[15232] == 15232 && 
b[15233] == 15233 && 
b[15234] == 15234 && 
b[15235] == 15235 && 
b[15236] == 15236 && 
b[15237] == 15237 && 
b[15238] == 15238 && 
b[15239] == 15239 && 
b[15240] == 15240 && 
b[15241] == 15241 && 
b[15242] == 15242 && 
b[15243] == 15243 && 
b[15244] == 15244 && 
b[15245] == 15245 && 
b[15246] == 15246 && 
b[15247] == 15247 && 
b[15248] == 15248 && 
b[15249] == 15249 && 
b[15250] == 15250 && 
b[15251] == 15251 && 
b[15252] == 15252 && 
b[15253] == 15253 && 
b[15254] == 15254 && 
b[15255] == 15255 && 
b[15256] == 15256 && 
b[15257] == 15257 && 
b[15258] == 15258 && 
b[15259] == 15259 && 
b[15260] == 15260 && 
b[15261] == 15261 && 
b[15262] == 15262 && 
b[15263] == 15263 && 
b[15264] == 15264 && 
b[15265] == 15265 && 
b[15266] == 15266 && 
b[15267] == 15267 && 
b[15268] == 15268 && 
b[15269] == 15269 && 
b[15270] == 15270 && 
b[15271] == 15271 && 
b[15272] == 15272 && 
b[15273] == 15273 && 
b[15274] == 15274 && 
b[15275] == 15275 && 
b[15276] == 15276 && 
b[15277] == 15277 && 
b[15278] == 15278 && 
b[15279] == 15279 && 
b[15280] == 15280 && 
b[15281] == 15281 && 
b[15282] == 15282 && 
b[15283] == 15283 && 
b[15284] == 15284 && 
b[15285] == 15285 && 
b[15286] == 15286 && 
b[15287] == 15287 && 
b[15288] == 15288 && 
b[15289] == 15289 && 
b[15290] == 15290 && 
b[15291] == 15291 && 
b[15292] == 15292 && 
b[15293] == 15293 && 
b[15294] == 15294 && 
b[15295] == 15295 && 
b[15296] == 15296 && 
b[15297] == 15297 && 
b[15298] == 15298 && 
b[15299] == 15299 && 
b[15300] == 15300 && 
b[15301] == 15301 && 
b[15302] == 15302 && 
b[15303] == 15303 && 
b[15304] == 15304 && 
b[15305] == 15305 && 
b[15306] == 15306 && 
b[15307] == 15307 && 
b[15308] == 15308 && 
b[15309] == 15309 && 
b[15310] == 15310 && 
b[15311] == 15311 && 
b[15312] == 15312 && 
b[15313] == 15313 && 
b[15314] == 15314 && 
b[15315] == 15315 && 
b[15316] == 15316 && 
b[15317] == 15317 && 
b[15318] == 15318 && 
b[15319] == 15319 && 
b[15320] == 15320 && 
b[15321] == 15321 && 
b[15322] == 15322 && 
b[15323] == 15323 && 
b[15324] == 15324 && 
b[15325] == 15325 && 
b[15326] == 15326 && 
b[15327] == 15327 && 
b[15328] == 15328 && 
b[15329] == 15329 && 
b[15330] == 15330 && 
b[15331] == 15331 && 
b[15332] == 15332 && 
b[15333] == 15333 && 
b[15334] == 15334 && 
b[15335] == 15335 && 
b[15336] == 15336 && 
b[15337] == 15337 && 
b[15338] == 15338 && 
b[15339] == 15339 && 
b[15340] == 15340 && 
b[15341] == 15341 && 
b[15342] == 15342 && 
b[15343] == 15343 && 
b[15344] == 15344 && 
b[15345] == 15345 && 
b[15346] == 15346 && 
b[15347] == 15347 && 
b[15348] == 15348 && 
b[15349] == 15349 && 
b[15350] == 15350 && 
b[15351] == 15351 && 
b[15352] == 15352 && 
b[15353] == 15353 && 
b[15354] == 15354 && 
b[15355] == 15355 && 
b[15356] == 15356 && 
b[15357] == 15357 && 
b[15358] == 15358 && 
b[15359] == 15359 && 
b[15360] == 15360 && 
b[15361] == 15361 && 
b[15362] == 15362 && 
b[15363] == 15363 && 
b[15364] == 15364 && 
b[15365] == 15365 && 
b[15366] == 15366 && 
b[15367] == 15367 && 
b[15368] == 15368 && 
b[15369] == 15369 && 
b[15370] == 15370 && 
b[15371] == 15371 && 
b[15372] == 15372 && 
b[15373] == 15373 && 
b[15374] == 15374 && 
b[15375] == 15375 && 
b[15376] == 15376 && 
b[15377] == 15377 && 
b[15378] == 15378 && 
b[15379] == 15379 && 
b[15380] == 15380 && 
b[15381] == 15381 && 
b[15382] == 15382 && 
b[15383] == 15383 && 
b[15384] == 15384 && 
b[15385] == 15385 && 
b[15386] == 15386 && 
b[15387] == 15387 && 
b[15388] == 15388 && 
b[15389] == 15389 && 
b[15390] == 15390 && 
b[15391] == 15391 && 
b[15392] == 15392 && 
b[15393] == 15393 && 
b[15394] == 15394 && 
b[15395] == 15395 && 
b[15396] == 15396 && 
b[15397] == 15397 && 
b[15398] == 15398 && 
b[15399] == 15399 && 
b[15400] == 15400 && 
b[15401] == 15401 && 
b[15402] == 15402 && 
b[15403] == 15403 && 
b[15404] == 15404 && 
b[15405] == 15405 && 
b[15406] == 15406 && 
b[15407] == 15407 && 
b[15408] == 15408 && 
b[15409] == 15409 && 
b[15410] == 15410 && 
b[15411] == 15411 && 
b[15412] == 15412 && 
b[15413] == 15413 && 
b[15414] == 15414 && 
b[15415] == 15415 && 
b[15416] == 15416 && 
b[15417] == 15417 && 
b[15418] == 15418 && 
b[15419] == 15419 && 
b[15420] == 15420 && 
b[15421] == 15421 && 
b[15422] == 15422 && 
b[15423] == 15423 && 
b[15424] == 15424 && 
b[15425] == 15425 && 
b[15426] == 15426 && 
b[15427] == 15427 && 
b[15428] == 15428 && 
b[15429] == 15429 && 
b[15430] == 15430 && 
b[15431] == 15431 && 
b[15432] == 15432 && 
b[15433] == 15433 && 
b[15434] == 15434 && 
b[15435] == 15435 && 
b[15436] == 15436 && 
b[15437] == 15437 && 
b[15438] == 15438 && 
b[15439] == 15439 && 
b[15440] == 15440 && 
b[15441] == 15441 && 
b[15442] == 15442 && 
b[15443] == 15443 && 
b[15444] == 15444 && 
b[15445] == 15445 && 
b[15446] == 15446 && 
b[15447] == 15447 && 
b[15448] == 15448 && 
b[15449] == 15449 && 
b[15450] == 15450 && 
b[15451] == 15451 && 
b[15452] == 15452 && 
b[15453] == 15453 && 
b[15454] == 15454 && 
b[15455] == 15455 && 
b[15456] == 15456 && 
b[15457] == 15457 && 
b[15458] == 15458 && 
b[15459] == 15459 && 
b[15460] == 15460 && 
b[15461] == 15461 && 
b[15462] == 15462 && 
b[15463] == 15463 && 
b[15464] == 15464 && 
b[15465] == 15465 && 
b[15466] == 15466 && 
b[15467] == 15467 && 
b[15468] == 15468 && 
b[15469] == 15469 && 
b[15470] == 15470 && 
b[15471] == 15471 && 
b[15472] == 15472 && 
b[15473] == 15473 && 
b[15474] == 15474 && 
b[15475] == 15475 && 
b[15476] == 15476 && 
b[15477] == 15477 && 
b[15478] == 15478 && 
b[15479] == 15479 && 
b[15480] == 15480 && 
b[15481] == 15481 && 
b[15482] == 15482 && 
b[15483] == 15483 && 
b[15484] == 15484 && 
b[15485] == 15485 && 
b[15486] == 15486 && 
b[15487] == 15487 && 
b[15488] == 15488 && 
b[15489] == 15489 && 
b[15490] == 15490 && 
b[15491] == 15491 && 
b[15492] == 15492 && 
b[15493] == 15493 && 
b[15494] == 15494 && 
b[15495] == 15495 && 
b[15496] == 15496 && 
b[15497] == 15497 && 
b[15498] == 15498 && 
b[15499] == 15499 && 
b[15500] == 15500 && 
b[15501] == 15501 && 
b[15502] == 15502 && 
b[15503] == 15503 && 
b[15504] == 15504 && 
b[15505] == 15505 && 
b[15506] == 15506 && 
b[15507] == 15507 && 
b[15508] == 15508 && 
b[15509] == 15509 && 
b[15510] == 15510 && 
b[15511] == 15511 && 
b[15512] == 15512 && 
b[15513] == 15513 && 
b[15514] == 15514 && 
b[15515] == 15515 && 
b[15516] == 15516 && 
b[15517] == 15517 && 
b[15518] == 15518 && 
b[15519] == 15519 && 
b[15520] == 15520 && 
b[15521] == 15521 && 
b[15522] == 15522 && 
b[15523] == 15523 && 
b[15524] == 15524 && 
b[15525] == 15525 && 
b[15526] == 15526 && 
b[15527] == 15527 && 
b[15528] == 15528 && 
b[15529] == 15529 && 
b[15530] == 15530 && 
b[15531] == 15531 && 
b[15532] == 15532 && 
b[15533] == 15533 && 
b[15534] == 15534 && 
b[15535] == 15535 && 
b[15536] == 15536 && 
b[15537] == 15537 && 
b[15538] == 15538 && 
b[15539] == 15539 && 
b[15540] == 15540 && 
b[15541] == 15541 && 
b[15542] == 15542 && 
b[15543] == 15543 && 
b[15544] == 15544 && 
b[15545] == 15545 && 
b[15546] == 15546 && 
b[15547] == 15547 && 
b[15548] == 15548 && 
b[15549] == 15549 && 
b[15550] == 15550 && 
b[15551] == 15551 && 
b[15552] == 15552 && 
b[15553] == 15553 && 
b[15554] == 15554 && 
b[15555] == 15555 && 
b[15556] == 15556 && 
b[15557] == 15557 && 
b[15558] == 15558 && 
b[15559] == 15559 && 
b[15560] == 15560 && 
b[15561] == 15561 && 
b[15562] == 15562 && 
b[15563] == 15563 && 
b[15564] == 15564 && 
b[15565] == 15565 && 
b[15566] == 15566 && 
b[15567] == 15567 && 
b[15568] == 15568 && 
b[15569] == 15569 && 
b[15570] == 15570 && 
b[15571] == 15571 && 
b[15572] == 15572 && 
b[15573] == 15573 && 
b[15574] == 15574 && 
b[15575] == 15575 && 
b[15576] == 15576 && 
b[15577] == 15577 && 
b[15578] == 15578 && 
b[15579] == 15579 && 
b[15580] == 15580 && 
b[15581] == 15581 && 
b[15582] == 15582 && 
b[15583] == 15583 && 
b[15584] == 15584 && 
b[15585] == 15585 && 
b[15586] == 15586 && 
b[15587] == 15587 && 
b[15588] == 15588 && 
b[15589] == 15589 && 
b[15590] == 15590 && 
b[15591] == 15591 && 
b[15592] == 15592 && 
b[15593] == 15593 && 
b[15594] == 15594 && 
b[15595] == 15595 && 
b[15596] == 15596 && 
b[15597] == 15597 && 
b[15598] == 15598 && 
b[15599] == 15599 && 
b[15600] == 15600 && 
b[15601] == 15601 && 
b[15602] == 15602 && 
b[15603] == 15603 && 
b[15604] == 15604 && 
b[15605] == 15605 && 
b[15606] == 15606 && 
b[15607] == 15607 && 
b[15608] == 15608 && 
b[15609] == 15609 && 
b[15610] == 15610 && 
b[15611] == 15611 && 
b[15612] == 15612 && 
b[15613] == 15613 && 
b[15614] == 15614 && 
b[15615] == 15615 && 
b[15616] == 15616 && 
b[15617] == 15617 && 
b[15618] == 15618 && 
b[15619] == 15619 && 
b[15620] == 15620 && 
b[15621] == 15621 && 
b[15622] == 15622 && 
b[15623] == 15623 && 
b[15624] == 15624 && 
b[15625] == 15625 && 
b[15626] == 15626 && 
b[15627] == 15627 && 
b[15628] == 15628 && 
b[15629] == 15629 && 
b[15630] == 15630 && 
b[15631] == 15631 && 
b[15632] == 15632 && 
b[15633] == 15633 && 
b[15634] == 15634 && 
b[15635] == 15635 && 
b[15636] == 15636 && 
b[15637] == 15637 && 
b[15638] == 15638 && 
b[15639] == 15639 && 
b[15640] == 15640 && 
b[15641] == 15641 && 
b[15642] == 15642 && 
b[15643] == 15643 && 
b[15644] == 15644 && 
b[15645] == 15645 && 
b[15646] == 15646 && 
b[15647] == 15647 && 
b[15648] == 15648 && 
b[15649] == 15649 && 
b[15650] == 15650 && 
b[15651] == 15651 && 
b[15652] == 15652 && 
b[15653] == 15653 && 
b[15654] == 15654 && 
b[15655] == 15655 && 
b[15656] == 15656 && 
b[15657] == 15657 && 
b[15658] == 15658 && 
b[15659] == 15659 && 
b[15660] == 15660 && 
b[15661] == 15661 && 
b[15662] == 15662 && 
b[15663] == 15663 && 
b[15664] == 15664 && 
b[15665] == 15665 && 
b[15666] == 15666 && 
b[15667] == 15667 && 
b[15668] == 15668 && 
b[15669] == 15669 && 
b[15670] == 15670 && 
b[15671] == 15671 && 
b[15672] == 15672 && 
b[15673] == 15673 && 
b[15674] == 15674 && 
b[15675] == 15675 && 
b[15676] == 15676 && 
b[15677] == 15677 && 
b[15678] == 15678 && 
b[15679] == 15679 && 
b[15680] == 15680 && 
b[15681] == 15681 && 
b[15682] == 15682 && 
b[15683] == 15683 && 
b[15684] == 15684 && 
b[15685] == 15685 && 
b[15686] == 15686 && 
b[15687] == 15687 && 
b[15688] == 15688 && 
b[15689] == 15689 && 
b[15690] == 15690 && 
b[15691] == 15691 && 
b[15692] == 15692 && 
b[15693] == 15693 && 
b[15694] == 15694 && 
b[15695] == 15695 && 
b[15696] == 15696 && 
b[15697] == 15697 && 
b[15698] == 15698 && 
b[15699] == 15699 && 
b[15700] == 15700 && 
b[15701] == 15701 && 
b[15702] == 15702 && 
b[15703] == 15703 && 
b[15704] == 15704 && 
b[15705] == 15705 && 
b[15706] == 15706 && 
b[15707] == 15707 && 
b[15708] == 15708 && 
b[15709] == 15709 && 
b[15710] == 15710 && 
b[15711] == 15711 && 
b[15712] == 15712 && 
b[15713] == 15713 && 
b[15714] == 15714 && 
b[15715] == 15715 && 
b[15716] == 15716 && 
b[15717] == 15717 && 
b[15718] == 15718 && 
b[15719] == 15719 && 
b[15720] == 15720 && 
b[15721] == 15721 && 
b[15722] == 15722 && 
b[15723] == 15723 && 
b[15724] == 15724 && 
b[15725] == 15725 && 
b[15726] == 15726 && 
b[15727] == 15727 && 
b[15728] == 15728 && 
b[15729] == 15729 && 
b[15730] == 15730 && 
b[15731] == 15731 && 
b[15732] == 15732 && 
b[15733] == 15733 && 
b[15734] == 15734 && 
b[15735] == 15735 && 
b[15736] == 15736 && 
b[15737] == 15737 && 
b[15738] == 15738 && 
b[15739] == 15739 && 
b[15740] == 15740 && 
b[15741] == 15741 && 
b[15742] == 15742 && 
b[15743] == 15743 && 
b[15744] == 15744 && 
b[15745] == 15745 && 
b[15746] == 15746 && 
b[15747] == 15747 && 
b[15748] == 15748 && 
b[15749] == 15749 && 
b[15750] == 15750 && 
b[15751] == 15751 && 
b[15752] == 15752 && 
b[15753] == 15753 && 
b[15754] == 15754 && 
b[15755] == 15755 && 
b[15756] == 15756 && 
b[15757] == 15757 && 
b[15758] == 15758 && 
b[15759] == 15759 && 
b[15760] == 15760 && 
b[15761] == 15761 && 
b[15762] == 15762 && 
b[15763] == 15763 && 
b[15764] == 15764 && 
b[15765] == 15765 && 
b[15766] == 15766 && 
b[15767] == 15767 && 
b[15768] == 15768 && 
b[15769] == 15769 && 
b[15770] == 15770 && 
b[15771] == 15771 && 
b[15772] == 15772 && 
b[15773] == 15773 && 
b[15774] == 15774 && 
b[15775] == 15775 && 
b[15776] == 15776 && 
b[15777] == 15777 && 
b[15778] == 15778 && 
b[15779] == 15779 && 
b[15780] == 15780 && 
b[15781] == 15781 && 
b[15782] == 15782 && 
b[15783] == 15783 && 
b[15784] == 15784 && 
b[15785] == 15785 && 
b[15786] == 15786 && 
b[15787] == 15787 && 
b[15788] == 15788 && 
b[15789] == 15789 && 
b[15790] == 15790 && 
b[15791] == 15791 && 
b[15792] == 15792 && 
b[15793] == 15793 && 
b[15794] == 15794 && 
b[15795] == 15795 && 
b[15796] == 15796 && 
b[15797] == 15797 && 
b[15798] == 15798 && 
b[15799] == 15799 && 
b[15800] == 15800 && 
b[15801] == 15801 && 
b[15802] == 15802 && 
b[15803] == 15803 && 
b[15804] == 15804 && 
b[15805] == 15805 && 
b[15806] == 15806 && 
b[15807] == 15807 && 
b[15808] == 15808 && 
b[15809] == 15809 && 
b[15810] == 15810 && 
b[15811] == 15811 && 
b[15812] == 15812 && 
b[15813] == 15813 && 
b[15814] == 15814 && 
b[15815] == 15815 && 
b[15816] == 15816 && 
b[15817] == 15817 && 
b[15818] == 15818 && 
b[15819] == 15819 && 
b[15820] == 15820 && 
b[15821] == 15821 && 
b[15822] == 15822 && 
b[15823] == 15823 && 
b[15824] == 15824 && 
b[15825] == 15825 && 
b[15826] == 15826 && 
b[15827] == 15827 && 
b[15828] == 15828 && 
b[15829] == 15829 && 
b[15830] == 15830 && 
b[15831] == 15831 && 
b[15832] == 15832 && 
b[15833] == 15833 && 
b[15834] == 15834 && 
b[15835] == 15835 && 
b[15836] == 15836 && 
b[15837] == 15837 && 
b[15838] == 15838 && 
b[15839] == 15839 && 
b[15840] == 15840 && 
b[15841] == 15841 && 
b[15842] == 15842 && 
b[15843] == 15843 && 
b[15844] == 15844 && 
b[15845] == 15845 && 
b[15846] == 15846 && 
b[15847] == 15847 && 
b[15848] == 15848 && 
b[15849] == 15849 && 
b[15850] == 15850 && 
b[15851] == 15851 && 
b[15852] == 15852 && 
b[15853] == 15853 && 
b[15854] == 15854 && 
b[15855] == 15855 && 
b[15856] == 15856 && 
b[15857] == 15857 && 
b[15858] == 15858 && 
b[15859] == 15859 && 
b[15860] == 15860 && 
b[15861] == 15861 && 
b[15862] == 15862 && 
b[15863] == 15863 && 
b[15864] == 15864 && 
b[15865] == 15865 && 
b[15866] == 15866 && 
b[15867] == 15867 && 
b[15868] == 15868 && 
b[15869] == 15869 && 
b[15870] == 15870 && 
b[15871] == 15871 && 
b[15872] == 15872 && 
b[15873] == 15873 && 
b[15874] == 15874 && 
b[15875] == 15875 && 
b[15876] == 15876 && 
b[15877] == 15877 && 
b[15878] == 15878 && 
b[15879] == 15879 && 
b[15880] == 15880 && 
b[15881] == 15881 && 
b[15882] == 15882 && 
b[15883] == 15883 && 
b[15884] == 15884 && 
b[15885] == 15885 && 
b[15886] == 15886 && 
b[15887] == 15887 && 
b[15888] == 15888 && 
b[15889] == 15889 && 
b[15890] == 15890 && 
b[15891] == 15891 && 
b[15892] == 15892 && 
b[15893] == 15893 && 
b[15894] == 15894 && 
b[15895] == 15895 && 
b[15896] == 15896 && 
b[15897] == 15897 && 
b[15898] == 15898 && 
b[15899] == 15899 && 
b[15900] == 15900 && 
b[15901] == 15901 && 
b[15902] == 15902 && 
b[15903] == 15903 && 
b[15904] == 15904 && 
b[15905] == 15905 && 
b[15906] == 15906 && 
b[15907] == 15907 && 
b[15908] == 15908 && 
b[15909] == 15909 && 
b[15910] == 15910 && 
b[15911] == 15911 && 
b[15912] == 15912 && 
b[15913] == 15913 && 
b[15914] == 15914 && 
b[15915] == 15915 && 
b[15916] == 15916 && 
b[15917] == 15917 && 
b[15918] == 15918 && 
b[15919] == 15919 && 
b[15920] == 15920 && 
b[15921] == 15921 && 
b[15922] == 15922 && 
b[15923] == 15923 && 
b[15924] == 15924 && 
b[15925] == 15925 && 
b[15926] == 15926 && 
b[15927] == 15927 && 
b[15928] == 15928 && 
b[15929] == 15929 && 
b[15930] == 15930 && 
b[15931] == 15931 && 
b[15932] == 15932 && 
b[15933] == 15933 && 
b[15934] == 15934 && 
b[15935] == 15935 && 
b[15936] == 15936 && 
b[15937] == 15937 && 
b[15938] == 15938 && 
b[15939] == 15939 && 
b[15940] == 15940 && 
b[15941] == 15941 && 
b[15942] == 15942 && 
b[15943] == 15943 && 
b[15944] == 15944 && 
b[15945] == 15945 && 
b[15946] == 15946 && 
b[15947] == 15947 && 
b[15948] == 15948 && 
b[15949] == 15949 && 
b[15950] == 15950 && 
b[15951] == 15951 && 
b[15952] == 15952 && 
b[15953] == 15953 && 
b[15954] == 15954 && 
b[15955] == 15955 && 
b[15956] == 15956 && 
b[15957] == 15957 && 
b[15958] == 15958 && 
b[15959] == 15959 && 
b[15960] == 15960 && 
b[15961] == 15961 && 
b[15962] == 15962 && 
b[15963] == 15963 && 
b[15964] == 15964 && 
b[15965] == 15965 && 
b[15966] == 15966 && 
b[15967] == 15967 && 
b[15968] == 15968 && 
b[15969] == 15969 && 
b[15970] == 15970 && 
b[15971] == 15971 && 
b[15972] == 15972 && 
b[15973] == 15973 && 
b[15974] == 15974 && 
b[15975] == 15975 && 
b[15976] == 15976 && 
b[15977] == 15977 && 
b[15978] == 15978 && 
b[15979] == 15979 && 
b[15980] == 15980 && 
b[15981] == 15981 && 
b[15982] == 15982 && 
b[15983] == 15983 && 
b[15984] == 15984 && 
b[15985] == 15985 && 
b[15986] == 15986 && 
b[15987] == 15987 && 
b[15988] == 15988 && 
b[15989] == 15989 && 
b[15990] == 15990 && 
b[15991] == 15991 && 
b[15992] == 15992 && 
b[15993] == 15993 && 
b[15994] == 15994 && 
b[15995] == 15995 && 
b[15996] == 15996 && 
b[15997] == 15997 && 
b[15998] == 15998 && 
b[15999] == 15999 && 
b[16000] == 16000 && 
b[16001] == 16001 && 
b[16002] == 16002 && 
b[16003] == 16003 && 
b[16004] == 16004 && 
b[16005] == 16005 && 
b[16006] == 16006 && 
b[16007] == 16007 && 
b[16008] == 16008 && 
b[16009] == 16009 && 
b[16010] == 16010 && 
b[16011] == 16011 && 
b[16012] == 16012 && 
b[16013] == 16013 && 
b[16014] == 16014 && 
b[16015] == 16015 && 
b[16016] == 16016 && 
b[16017] == 16017 && 
b[16018] == 16018 && 
b[16019] == 16019 && 
b[16020] == 16020 && 
b[16021] == 16021 && 
b[16022] == 16022 && 
b[16023] == 16023 && 
b[16024] == 16024 && 
b[16025] == 16025 && 
b[16026] == 16026 && 
b[16027] == 16027 && 
b[16028] == 16028 && 
b[16029] == 16029 && 
b[16030] == 16030 && 
b[16031] == 16031 && 
b[16032] == 16032 && 
b[16033] == 16033 && 
b[16034] == 16034 && 
b[16035] == 16035 && 
b[16036] == 16036 && 
b[16037] == 16037 && 
b[16038] == 16038 && 
b[16039] == 16039 && 
b[16040] == 16040 && 
b[16041] == 16041 && 
b[16042] == 16042 && 
b[16043] == 16043 && 
b[16044] == 16044 && 
b[16045] == 16045 && 
b[16046] == 16046 && 
b[16047] == 16047 && 
b[16048] == 16048 && 
b[16049] == 16049 && 
b[16050] == 16050 && 
b[16051] == 16051 && 
b[16052] == 16052 && 
b[16053] == 16053 && 
b[16054] == 16054 && 
b[16055] == 16055 && 
b[16056] == 16056 && 
b[16057] == 16057 && 
b[16058] == 16058 && 
b[16059] == 16059 && 
b[16060] == 16060 && 
b[16061] == 16061 && 
b[16062] == 16062 && 
b[16063] == 16063 && 
b[16064] == 16064 && 
b[16065] == 16065 && 
b[16066] == 16066 && 
b[16067] == 16067 && 
b[16068] == 16068 && 
b[16069] == 16069 && 
b[16070] == 16070 && 
b[16071] == 16071 && 
b[16072] == 16072 && 
b[16073] == 16073 && 
b[16074] == 16074 && 
b[16075] == 16075 && 
b[16076] == 16076 && 
b[16077] == 16077 && 
b[16078] == 16078 && 
b[16079] == 16079 && 
b[16080] == 16080 && 
b[16081] == 16081 && 
b[16082] == 16082 && 
b[16083] == 16083 && 
b[16084] == 16084 && 
b[16085] == 16085 && 
b[16086] == 16086 && 
b[16087] == 16087 && 
b[16088] == 16088 && 
b[16089] == 16089 && 
b[16090] == 16090 && 
b[16091] == 16091 && 
b[16092] == 16092 && 
b[16093] == 16093 && 
b[16094] == 16094 && 
b[16095] == 16095 && 
b[16096] == 16096 && 
b[16097] == 16097 && 
b[16098] == 16098 && 
b[16099] == 16099 && 
b[16100] == 16100 && 
b[16101] == 16101 && 
b[16102] == 16102 && 
b[16103] == 16103 && 
b[16104] == 16104 && 
b[16105] == 16105 && 
b[16106] == 16106 && 
b[16107] == 16107 && 
b[16108] == 16108 && 
b[16109] == 16109 && 
b[16110] == 16110 && 
b[16111] == 16111 && 
b[16112] == 16112 && 
b[16113] == 16113 && 
b[16114] == 16114 && 
b[16115] == 16115 && 
b[16116] == 16116 && 
b[16117] == 16117 && 
b[16118] == 16118 && 
b[16119] == 16119 && 
b[16120] == 16120 && 
b[16121] == 16121 && 
b[16122] == 16122 && 
b[16123] == 16123 && 
b[16124] == 16124 && 
b[16125] == 16125 && 
b[16126] == 16126 && 
b[16127] == 16127 && 
b[16128] == 16128 && 
b[16129] == 16129 && 
b[16130] == 16130 && 
b[16131] == 16131 && 
b[16132] == 16132 && 
b[16133] == 16133 && 
b[16134] == 16134 && 
b[16135] == 16135 && 
b[16136] == 16136 && 
b[16137] == 16137 && 
b[16138] == 16138 && 
b[16139] == 16139 && 
b[16140] == 16140 && 
b[16141] == 16141 && 
b[16142] == 16142 && 
b[16143] == 16143 && 
b[16144] == 16144 && 
b[16145] == 16145 && 
b[16146] == 16146 && 
b[16147] == 16147 && 
b[16148] == 16148 && 
b[16149] == 16149 && 
b[16150] == 16150 && 
b[16151] == 16151 && 
b[16152] == 16152 && 
b[16153] == 16153 && 
b[16154] == 16154 && 
b[16155] == 16155 && 
b[16156] == 16156 && 
b[16157] == 16157 && 
b[16158] == 16158 && 
b[16159] == 16159 && 
b[16160] == 16160 && 
b[16161] == 16161 && 
b[16162] == 16162 && 
b[16163] == 16163 && 
b[16164] == 16164 && 
b[16165] == 16165 && 
b[16166] == 16166 && 
b[16167] == 16167 && 
b[16168] == 16168 && 
b[16169] == 16169 && 
b[16170] == 16170 && 
b[16171] == 16171 && 
b[16172] == 16172 && 
b[16173] == 16173 && 
b[16174] == 16174 && 
b[16175] == 16175 && 
b[16176] == 16176 && 
b[16177] == 16177 && 
b[16178] == 16178 && 
b[16179] == 16179 && 
b[16180] == 16180 && 
b[16181] == 16181 && 
b[16182] == 16182 && 
b[16183] == 16183 && 
b[16184] == 16184 && 
b[16185] == 16185 && 
b[16186] == 16186 && 
b[16187] == 16187 && 
b[16188] == 16188 && 
b[16189] == 16189 && 
b[16190] == 16190 && 
b[16191] == 16191 && 
b[16192] == 16192 && 
b[16193] == 16193 && 
b[16194] == 16194 && 
b[16195] == 16195 && 
b[16196] == 16196 && 
b[16197] == 16197 && 
b[16198] == 16198 && 
b[16199] == 16199 && 
b[16200] == 16200 && 
b[16201] == 16201 && 
b[16202] == 16202 && 
b[16203] == 16203 && 
b[16204] == 16204 && 
b[16205] == 16205 && 
b[16206] == 16206 && 
b[16207] == 16207 && 
b[16208] == 16208 && 
b[16209] == 16209 && 
b[16210] == 16210 && 
b[16211] == 16211 && 
b[16212] == 16212 && 
b[16213] == 16213 && 
b[16214] == 16214 && 
b[16215] == 16215 && 
b[16216] == 16216 && 
b[16217] == 16217 && 
b[16218] == 16218 && 
b[16219] == 16219 && 
b[16220] == 16220 && 
b[16221] == 16221 && 
b[16222] == 16222 && 
b[16223] == 16223 && 
b[16224] == 16224 && 
b[16225] == 16225 && 
b[16226] == 16226 && 
b[16227] == 16227 && 
b[16228] == 16228 && 
b[16229] == 16229 && 
b[16230] == 16230 && 
b[16231] == 16231 && 
b[16232] == 16232 && 
b[16233] == 16233 && 
b[16234] == 16234 && 
b[16235] == 16235 && 
b[16236] == 16236 && 
b[16237] == 16237 && 
b[16238] == 16238 && 
b[16239] == 16239 && 
b[16240] == 16240 && 
b[16241] == 16241 && 
b[16242] == 16242 && 
b[16243] == 16243 && 
b[16244] == 16244 && 
b[16245] == 16245 && 
b[16246] == 16246 && 
b[16247] == 16247 && 
b[16248] == 16248 && 
b[16249] == 16249 && 
b[16250] == 16250 && 
b[16251] == 16251 && 
b[16252] == 16252 && 
b[16253] == 16253 && 
b[16254] == 16254 && 
b[16255] == 16255 && 
b[16256] == 16256 && 
b[16257] == 16257 && 
b[16258] == 16258 && 
b[16259] == 16259 && 
b[16260] == 16260 && 
b[16261] == 16261 && 
b[16262] == 16262 && 
b[16263] == 16263 && 
b[16264] == 16264 && 
b[16265] == 16265 && 
b[16266] == 16266 && 
b[16267] == 16267 && 
b[16268] == 16268 && 
b[16269] == 16269 && 
b[16270] == 16270 && 
b[16271] == 16271 && 
b[16272] == 16272 && 
b[16273] == 16273 && 
b[16274] == 16274 && 
b[16275] == 16275 && 
b[16276] == 16276 && 
b[16277] == 16277 && 
b[16278] == 16278 && 
b[16279] == 16279 && 
b[16280] == 16280 && 
b[16281] == 16281 && 
b[16282] == 16282 && 
b[16283] == 16283 && 
b[16284] == 16284 && 
b[16285] == 16285 && 
b[16286] == 16286 && 
b[16287] == 16287 && 
b[16288] == 16288 && 
b[16289] == 16289 && 
b[16290] == 16290 && 
b[16291] == 16291 && 
b[16292] == 16292 && 
b[16293] == 16293 && 
b[16294] == 16294 && 
b[16295] == 16295 && 
b[16296] == 16296 && 
b[16297] == 16297 && 
b[16298] == 16298 && 
b[16299] == 16299 && 
b[16300] == 16300 && 
b[16301] == 16301 && 
b[16302] == 16302 && 
b[16303] == 16303 && 
b[16304] == 16304 && 
b[16305] == 16305 && 
b[16306] == 16306 && 
b[16307] == 16307 && 
b[16308] == 16308 && 
b[16309] == 16309 && 
b[16310] == 16310 && 
b[16311] == 16311 && 
b[16312] == 16312 && 
b[16313] == 16313 && 
b[16314] == 16314 && 
b[16315] == 16315 && 
b[16316] == 16316 && 
b[16317] == 16317 && 
b[16318] == 16318 && 
b[16319] == 16319 && 
b[16320] == 16320 && 
b[16321] == 16321 && 
b[16322] == 16322 && 
b[16323] == 16323 && 
b[16324] == 16324 && 
b[16325] == 16325 && 
b[16326] == 16326 && 
b[16327] == 16327 && 
b[16328] == 16328 && 
b[16329] == 16329 && 
b[16330] == 16330 && 
b[16331] == 16331 && 
b[16332] == 16332 && 
b[16333] == 16333 && 
b[16334] == 16334 && 
b[16335] == 16335 && 
b[16336] == 16336 && 
b[16337] == 16337 && 
b[16338] == 16338 && 
b[16339] == 16339 && 
b[16340] == 16340 && 
b[16341] == 16341 && 
b[16342] == 16342 && 
b[16343] == 16343 && 
b[16344] == 16344 && 
b[16345] == 16345 && 
b[16346] == 16346 && 
b[16347] == 16347 && 
b[16348] == 16348 && 
b[16349] == 16349 && 
b[16350] == 16350 && 
b[16351] == 16351 && 
b[16352] == 16352 && 
b[16353] == 16353 && 
b[16354] == 16354 && 
b[16355] == 16355 && 
b[16356] == 16356 && 
b[16357] == 16357 && 
b[16358] == 16358 && 
b[16359] == 16359 && 
b[16360] == 16360 && 
b[16361] == 16361 && 
b[16362] == 16362 && 
b[16363] == 16363 && 
b[16364] == 16364 && 
b[16365] == 16365 && 
b[16366] == 16366 && 
b[16367] == 16367 && 
b[16368] == 16368 && 
b[16369] == 16369 && 
b[16370] == 16370 && 
b[16371] == 16371 && 
b[16372] == 16372 && 
b[16373] == 16373 && 
b[16374] == 16374 && 
b[16375] == 16375 && 
b[16376] == 16376 && 
b[16377] == 16377 && 
b[16378] == 16378 && 
b[16379] == 16379 && 
b[16380] == 16380 && 
b[16381] == 16381 && 
b[16382] == 16382 && 
b[16383] == 16383 && 
b[16384] == 16384 && 
b[16385] == 16385 && 
b[16386] == 16386 && 
b[16387] == 16387 && 
b[16388] == 16388 && 
b[16389] == 16389 && 
b[16390] == 16390 && 
b[16391] == 16391 && 
b[16392] == 16392 && 
b[16393] == 16393 && 
b[16394] == 16394 && 
b[16395] == 16395 && 
b[16396] == 16396 && 
b[16397] == 16397 && 
b[16398] == 16398 && 
b[16399] == 16399 && 
b[16400] == 16400 && 
b[16401] == 16401 && 
b[16402] == 16402 && 
b[16403] == 16403 && 
b[16404] == 16404 && 
b[16405] == 16405 && 
b[16406] == 16406 && 
b[16407] == 16407 && 
b[16408] == 16408 && 
b[16409] == 16409 && 
b[16410] == 16410 && 
b[16411] == 16411 && 
b[16412] == 16412 && 
b[16413] == 16413 && 
b[16414] == 16414 && 
b[16415] == 16415 && 
b[16416] == 16416 && 
b[16417] == 16417 && 
b[16418] == 16418 && 
b[16419] == 16419 && 
b[16420] == 16420 && 
b[16421] == 16421 && 
b[16422] == 16422 && 
b[16423] == 16423 && 
b[16424] == 16424 && 
b[16425] == 16425 && 
b[16426] == 16426 && 
b[16427] == 16427 && 
b[16428] == 16428 && 
b[16429] == 16429 && 
b[16430] == 16430 && 
b[16431] == 16431 && 
b[16432] == 16432 && 
b[16433] == 16433 && 
b[16434] == 16434 && 
b[16435] == 16435 && 
b[16436] == 16436 && 
b[16437] == 16437 && 
b[16438] == 16438 && 
b[16439] == 16439 && 
b[16440] == 16440 && 
b[16441] == 16441 && 
b[16442] == 16442 && 
b[16443] == 16443 && 
b[16444] == 16444 && 
b[16445] == 16445 && 
b[16446] == 16446 && 
b[16447] == 16447 && 
b[16448] == 16448 && 
b[16449] == 16449 && 
b[16450] == 16450 && 
b[16451] == 16451 && 
b[16452] == 16452 && 
b[16453] == 16453 && 
b[16454] == 16454 && 
b[16455] == 16455 && 
b[16456] == 16456 && 
b[16457] == 16457 && 
b[16458] == 16458 && 
b[16459] == 16459 && 
b[16460] == 16460 && 
b[16461] == 16461 && 
b[16462] == 16462 && 
b[16463] == 16463 && 
b[16464] == 16464 && 
b[16465] == 16465 && 
b[16466] == 16466 && 
b[16467] == 16467 && 
b[16468] == 16468 && 
b[16469] == 16469 && 
b[16470] == 16470 && 
b[16471] == 16471 && 
b[16472] == 16472 && 
b[16473] == 16473 && 
b[16474] == 16474 && 
b[16475] == 16475 && 
b[16476] == 16476 && 
b[16477] == 16477 && 
b[16478] == 16478 && 
b[16479] == 16479 && 
b[16480] == 16480 && 
b[16481] == 16481 && 
b[16482] == 16482 && 
b[16483] == 16483 && 
b[16484] == 16484 && 
b[16485] == 16485 && 
b[16486] == 16486 && 
b[16487] == 16487 && 
b[16488] == 16488 && 
b[16489] == 16489 && 
b[16490] == 16490 && 
b[16491] == 16491 && 
b[16492] == 16492 && 
b[16493] == 16493 && 
b[16494] == 16494 && 
b[16495] == 16495 && 
b[16496] == 16496 && 
b[16497] == 16497 && 
b[16498] == 16498 && 
b[16499] == 16499 && 
b[16500] == 16500 && 
b[16501] == 16501 && 
b[16502] == 16502 && 
b[16503] == 16503 && 
b[16504] == 16504 && 
b[16505] == 16505 && 
b[16506] == 16506 && 
b[16507] == 16507 && 
b[16508] == 16508 && 
b[16509] == 16509 && 
b[16510] == 16510 && 
b[16511] == 16511 && 
b[16512] == 16512 && 
b[16513] == 16513 && 
b[16514] == 16514 && 
b[16515] == 16515 && 
b[16516] == 16516 && 
b[16517] == 16517 && 
b[16518] == 16518 && 
b[16519] == 16519 && 
b[16520] == 16520 && 
b[16521] == 16521 && 
b[16522] == 16522 && 
b[16523] == 16523 && 
b[16524] == 16524 && 
b[16525] == 16525 && 
b[16526] == 16526 && 
b[16527] == 16527 && 
b[16528] == 16528 && 
b[16529] == 16529 && 
b[16530] == 16530 && 
b[16531] == 16531 && 
b[16532] == 16532 && 
b[16533] == 16533 && 
b[16534] == 16534 && 
b[16535] == 16535 && 
b[16536] == 16536 && 
b[16537] == 16537 && 
b[16538] == 16538 && 
b[16539] == 16539 && 
b[16540] == 16540 && 
b[16541] == 16541 && 
b[16542] == 16542 && 
b[16543] == 16543 && 
b[16544] == 16544 && 
b[16545] == 16545 && 
b[16546] == 16546 && 
b[16547] == 16547 && 
b[16548] == 16548 && 
b[16549] == 16549 && 
b[16550] == 16550 && 
b[16551] == 16551 && 
b[16552] == 16552 && 
b[16553] == 16553 && 
b[16554] == 16554 && 
b[16555] == 16555 && 
b[16556] == 16556 && 
b[16557] == 16557 && 
b[16558] == 16558 && 
b[16559] == 16559 && 
b[16560] == 16560 && 
b[16561] == 16561 && 
b[16562] == 16562 && 
b[16563] == 16563 && 
b[16564] == 16564 && 
b[16565] == 16565 && 
b[16566] == 16566 && 
b[16567] == 16567 && 
b[16568] == 16568 && 
b[16569] == 16569 && 
b[16570] == 16570 && 
b[16571] == 16571 && 
b[16572] == 16572 && 
b[16573] == 16573 && 
b[16574] == 16574 && 
b[16575] == 16575 && 
b[16576] == 16576 && 
b[16577] == 16577 && 
b[16578] == 16578 && 
b[16579] == 16579 && 
b[16580] == 16580 && 
b[16581] == 16581 && 
b[16582] == 16582 && 
b[16583] == 16583 && 
b[16584] == 16584 && 
b[16585] == 16585 && 
b[16586] == 16586 && 
b[16587] == 16587 && 
b[16588] == 16588 && 
b[16589] == 16589 && 
b[16590] == 16590 && 
b[16591] == 16591 && 
b[16592] == 16592 && 
b[16593] == 16593 && 
b[16594] == 16594 && 
b[16595] == 16595 && 
b[16596] == 16596 && 
b[16597] == 16597 && 
b[16598] == 16598 && 
b[16599] == 16599 && 
b[16600] == 16600 && 
b[16601] == 16601 && 
b[16602] == 16602 && 
b[16603] == 16603 && 
b[16604] == 16604 && 
b[16605] == 16605 && 
b[16606] == 16606 && 
b[16607] == 16607 && 
b[16608] == 16608 && 
b[16609] == 16609 && 
b[16610] == 16610 && 
b[16611] == 16611 && 
b[16612] == 16612 && 
b[16613] == 16613 && 
b[16614] == 16614 && 
b[16615] == 16615 && 
b[16616] == 16616 && 
b[16617] == 16617 && 
b[16618] == 16618 && 
b[16619] == 16619 && 
b[16620] == 16620 && 
b[16621] == 16621 && 
b[16622] == 16622 && 
b[16623] == 16623 && 
b[16624] == 16624 && 
b[16625] == 16625 && 
b[16626] == 16626 && 
b[16627] == 16627 && 
b[16628] == 16628 && 
b[16629] == 16629 && 
b[16630] == 16630 && 
b[16631] == 16631 && 
b[16632] == 16632 && 
b[16633] == 16633 && 
b[16634] == 16634 && 
b[16635] == 16635 && 
b[16636] == 16636 && 
b[16637] == 16637 && 
b[16638] == 16638 && 
b[16639] == 16639 && 
b[16640] == 16640 && 
b[16641] == 16641 && 
b[16642] == 16642 && 
b[16643] == 16643 && 
b[16644] == 16644 && 
b[16645] == 16645 && 
b[16646] == 16646 && 
b[16647] == 16647 && 
b[16648] == 16648 && 
b[16649] == 16649 && 
b[16650] == 16650 && 
b[16651] == 16651 && 
b[16652] == 16652 && 
b[16653] == 16653 && 
b[16654] == 16654 && 
b[16655] == 16655 && 
b[16656] == 16656 && 
b[16657] == 16657 && 
b[16658] == 16658 && 
b[16659] == 16659 && 
b[16660] == 16660 && 
b[16661] == 16661 && 
b[16662] == 16662 && 
b[16663] == 16663 && 
b[16664] == 16664 && 
b[16665] == 16665 && 
b[16666] == 16666 && 
b[16667] == 16667 && 
b[16668] == 16668 && 
b[16669] == 16669 && 
b[16670] == 16670 && 
b[16671] == 16671 && 
b[16672] == 16672 && 
b[16673] == 16673 && 
b[16674] == 16674 && 
b[16675] == 16675 && 
b[16676] == 16676 && 
b[16677] == 16677 && 
b[16678] == 16678 && 
b[16679] == 16679 && 
b[16680] == 16680 && 
b[16681] == 16681 && 
b[16682] == 16682 && 
b[16683] == 16683 && 
b[16684] == 16684 && 
b[16685] == 16685 && 
b[16686] == 16686 && 
b[16687] == 16687 && 
b[16688] == 16688 && 
b[16689] == 16689 && 
b[16690] == 16690 && 
b[16691] == 16691 && 
b[16692] == 16692 && 
b[16693] == 16693 && 
b[16694] == 16694 && 
b[16695] == 16695 && 
b[16696] == 16696 && 
b[16697] == 16697 && 
b[16698] == 16698 && 
b[16699] == 16699 && 
b[16700] == 16700 && 
b[16701] == 16701 && 
b[16702] == 16702 && 
b[16703] == 16703 && 
b[16704] == 16704 && 
b[16705] == 16705 && 
b[16706] == 16706 && 
b[16707] == 16707 && 
b[16708] == 16708 && 
b[16709] == 16709 && 
b[16710] == 16710 && 
b[16711] == 16711 && 
b[16712] == 16712 && 
b[16713] == 16713 && 
b[16714] == 16714 && 
b[16715] == 16715 && 
b[16716] == 16716 && 
b[16717] == 16717 && 
b[16718] == 16718 && 
b[16719] == 16719 && 
b[16720] == 16720 && 
b[16721] == 16721 && 
b[16722] == 16722 && 
b[16723] == 16723 && 
b[16724] == 16724 && 
b[16725] == 16725 && 
b[16726] == 16726 && 
b[16727] == 16727 && 
b[16728] == 16728 && 
b[16729] == 16729 && 
b[16730] == 16730 && 
b[16731] == 16731 && 
b[16732] == 16732 && 
b[16733] == 16733 && 
b[16734] == 16734 && 
b[16735] == 16735 && 
b[16736] == 16736 && 
b[16737] == 16737 && 
b[16738] == 16738 && 
b[16739] == 16739 && 
b[16740] == 16740 && 
b[16741] == 16741 && 
b[16742] == 16742 && 
b[16743] == 16743 && 
b[16744] == 16744 && 
b[16745] == 16745 && 
b[16746] == 16746 && 
b[16747] == 16747 && 
b[16748] == 16748 && 
b[16749] == 16749 && 
b[16750] == 16750 && 
b[16751] == 16751 && 
b[16752] == 16752 && 
b[16753] == 16753 && 
b[16754] == 16754 && 
b[16755] == 16755 && 
b[16756] == 16756 && 
b[16757] == 16757 && 
b[16758] == 16758 && 
b[16759] == 16759 && 
b[16760] == 16760 && 
b[16761] == 16761 && 
b[16762] == 16762 && 
b[16763] == 16763 && 
b[16764] == 16764 && 
b[16765] == 16765 && 
b[16766] == 16766 && 
b[16767] == 16767 && 
b[16768] == 16768 && 
b[16769] == 16769 && 
b[16770] == 16770 && 
b[16771] == 16771 && 
b[16772] == 16772 && 
b[16773] == 16773 && 
b[16774] == 16774 && 
b[16775] == 16775 && 
b[16776] == 16776 && 
b[16777] == 16777 && 
b[16778] == 16778 && 
b[16779] == 16779 && 
b[16780] == 16780 && 
b[16781] == 16781 && 
b[16782] == 16782 && 
b[16783] == 16783 && 
b[16784] == 16784 && 
b[16785] == 16785 && 
b[16786] == 16786 && 
b[16787] == 16787 && 
b[16788] == 16788 && 
b[16789] == 16789 && 
b[16790] == 16790 && 
b[16791] == 16791 && 
b[16792] == 16792 && 
b[16793] == 16793 && 
b[16794] == 16794 && 
b[16795] == 16795 && 
b[16796] == 16796 && 
b[16797] == 16797 && 
b[16798] == 16798 && 
b[16799] == 16799 && 
b[16800] == 16800 && 
b[16801] == 16801 && 
b[16802] == 16802 && 
b[16803] == 16803 && 
b[16804] == 16804 && 
b[16805] == 16805 && 
b[16806] == 16806 && 
b[16807] == 16807 && 
b[16808] == 16808 && 
b[16809] == 16809 && 
b[16810] == 16810 && 
b[16811] == 16811 && 
b[16812] == 16812 && 
b[16813] == 16813 && 
b[16814] == 16814 && 
b[16815] == 16815 && 
b[16816] == 16816 && 
b[16817] == 16817 && 
b[16818] == 16818 && 
b[16819] == 16819 && 
b[16820] == 16820 && 
b[16821] == 16821 && 
b[16822] == 16822 && 
b[16823] == 16823 && 
b[16824] == 16824 && 
b[16825] == 16825 && 
b[16826] == 16826 && 
b[16827] == 16827 && 
b[16828] == 16828 && 
b[16829] == 16829 && 
b[16830] == 16830 && 
b[16831] == 16831 && 
b[16832] == 16832 && 
b[16833] == 16833 && 
b[16834] == 16834 && 
b[16835] == 16835 && 
b[16836] == 16836 && 
b[16837] == 16837 && 
b[16838] == 16838 && 
b[16839] == 16839 && 
b[16840] == 16840 && 
b[16841] == 16841 && 
b[16842] == 16842 && 
b[16843] == 16843 && 
b[16844] == 16844 && 
b[16845] == 16845 && 
b[16846] == 16846 && 
b[16847] == 16847 && 
b[16848] == 16848 && 
b[16849] == 16849 && 
b[16850] == 16850 && 
b[16851] == 16851 && 
b[16852] == 16852 && 
b[16853] == 16853 && 
b[16854] == 16854 && 
b[16855] == 16855 && 
b[16856] == 16856 && 
b[16857] == 16857 && 
b[16858] == 16858 && 
b[16859] == 16859 && 
b[16860] == 16860 && 
b[16861] == 16861 && 
b[16862] == 16862 && 
b[16863] == 16863 && 
b[16864] == 16864 && 
b[16865] == 16865 && 
b[16866] == 16866 && 
b[16867] == 16867 && 
b[16868] == 16868 && 
b[16869] == 16869 && 
b[16870] == 16870 && 
b[16871] == 16871 && 
b[16872] == 16872 && 
b[16873] == 16873 && 
b[16874] == 16874 && 
b[16875] == 16875 && 
b[16876] == 16876 && 
b[16877] == 16877 && 
b[16878] == 16878 && 
b[16879] == 16879 && 
b[16880] == 16880 && 
b[16881] == 16881 && 
b[16882] == 16882 && 
b[16883] == 16883 && 
b[16884] == 16884 && 
b[16885] == 16885 && 
b[16886] == 16886 && 
b[16887] == 16887 && 
b[16888] == 16888 && 
b[16889] == 16889 && 
b[16890] == 16890 && 
b[16891] == 16891 && 
b[16892] == 16892 && 
b[16893] == 16893 && 
b[16894] == 16894 && 
b[16895] == 16895 && 
b[16896] == 16896 && 
b[16897] == 16897 && 
b[16898] == 16898 && 
b[16899] == 16899 && 
b[16900] == 16900 && 
b[16901] == 16901 && 
b[16902] == 16902 && 
b[16903] == 16903 && 
b[16904] == 16904 && 
b[16905] == 16905 && 
b[16906] == 16906 && 
b[16907] == 16907 && 
b[16908] == 16908 && 
b[16909] == 16909 && 
b[16910] == 16910 && 
b[16911] == 16911 && 
b[16912] == 16912 && 
b[16913] == 16913 && 
b[16914] == 16914 && 
b[16915] == 16915 && 
b[16916] == 16916 && 
b[16917] == 16917 && 
b[16918] == 16918 && 
b[16919] == 16919 && 
b[16920] == 16920 && 
b[16921] == 16921 && 
b[16922] == 16922 && 
b[16923] == 16923 && 
b[16924] == 16924 && 
b[16925] == 16925 && 
b[16926] == 16926 && 
b[16927] == 16927 && 
b[16928] == 16928 && 
b[16929] == 16929 && 
b[16930] == 16930 && 
b[16931] == 16931 && 
b[16932] == 16932 && 
b[16933] == 16933 && 
b[16934] == 16934 && 
b[16935] == 16935 && 
b[16936] == 16936 && 
b[16937] == 16937 && 
b[16938] == 16938 && 
b[16939] == 16939 && 
b[16940] == 16940 && 
b[16941] == 16941 && 
b[16942] == 16942 && 
b[16943] == 16943 && 
b[16944] == 16944 && 
b[16945] == 16945 && 
b[16946] == 16946 && 
b[16947] == 16947 && 
b[16948] == 16948 && 
b[16949] == 16949 && 
b[16950] == 16950 && 
b[16951] == 16951 && 
b[16952] == 16952 && 
b[16953] == 16953 && 
b[16954] == 16954 && 
b[16955] == 16955 && 
b[16956] == 16956 && 
b[16957] == 16957 && 
b[16958] == 16958 && 
b[16959] == 16959 && 
b[16960] == 16960 && 
b[16961] == 16961 && 
b[16962] == 16962 && 
b[16963] == 16963 && 
b[16964] == 16964 && 
b[16965] == 16965 && 
b[16966] == 16966 && 
b[16967] == 16967 && 
b[16968] == 16968 && 
b[16969] == 16969 && 
b[16970] == 16970 && 
b[16971] == 16971 && 
b[16972] == 16972 && 
b[16973] == 16973 && 
b[16974] == 16974 && 
b[16975] == 16975 && 
b[16976] == 16976 && 
b[16977] == 16977 && 
b[16978] == 16978 && 
b[16979] == 16979 && 
b[16980] == 16980 && 
b[16981] == 16981 && 
b[16982] == 16982 && 
b[16983] == 16983 && 
b[16984] == 16984 && 
b[16985] == 16985 && 
b[16986] == 16986 && 
b[16987] == 16987 && 
b[16988] == 16988 && 
b[16989] == 16989 && 
b[16990] == 16990 && 
b[16991] == 16991 && 
b[16992] == 16992 && 
b[16993] == 16993 && 
b[16994] == 16994 && 
b[16995] == 16995 && 
b[16996] == 16996 && 
b[16997] == 16997 && 
b[16998] == 16998 && 
b[16999] == 16999 && 
b[17000] == 17000 && 
b[17001] == 17001 && 
b[17002] == 17002 && 
b[17003] == 17003 && 
b[17004] == 17004 && 
b[17005] == 17005 && 
b[17006] == 17006 && 
b[17007] == 17007 && 
b[17008] == 17008 && 
b[17009] == 17009 && 
b[17010] == 17010 && 
b[17011] == 17011 && 
b[17012] == 17012 && 
b[17013] == 17013 && 
b[17014] == 17014 && 
b[17015] == 17015 && 
b[17016] == 17016 && 
b[17017] == 17017 && 
b[17018] == 17018 && 
b[17019] == 17019 && 
b[17020] == 17020 && 
b[17021] == 17021 && 
b[17022] == 17022 && 
b[17023] == 17023 && 
b[17024] == 17024 && 
b[17025] == 17025 && 
b[17026] == 17026 && 
b[17027] == 17027 && 
b[17028] == 17028 && 
b[17029] == 17029 && 
b[17030] == 17030 && 
b[17031] == 17031 && 
b[17032] == 17032 && 
b[17033] == 17033 && 
b[17034] == 17034 && 
b[17035] == 17035 && 
b[17036] == 17036 && 
b[17037] == 17037 && 
b[17038] == 17038 && 
b[17039] == 17039 && 
b[17040] == 17040 && 
b[17041] == 17041 && 
b[17042] == 17042 && 
b[17043] == 17043 && 
b[17044] == 17044 && 
b[17045] == 17045 && 
b[17046] == 17046 && 
b[17047] == 17047 && 
b[17048] == 17048 && 
b[17049] == 17049 && 
b[17050] == 17050 && 
b[17051] == 17051 && 
b[17052] == 17052 && 
b[17053] == 17053 && 
b[17054] == 17054 && 
b[17055] == 17055 && 
b[17056] == 17056 && 
b[17057] == 17057 && 
b[17058] == 17058 && 
b[17059] == 17059 && 
b[17060] == 17060 && 
b[17061] == 17061 && 
b[17062] == 17062 && 
b[17063] == 17063 && 
b[17064] == 17064 && 
b[17065] == 17065 && 
b[17066] == 17066 && 
b[17067] == 17067 && 
b[17068] == 17068 && 
b[17069] == 17069 && 
b[17070] == 17070 && 
b[17071] == 17071 && 
b[17072] == 17072 && 
b[17073] == 17073 && 
b[17074] == 17074 && 
b[17075] == 17075 && 
b[17076] == 17076 && 
b[17077] == 17077 && 
b[17078] == 17078 && 
b[17079] == 17079 && 
b[17080] == 17080 && 
b[17081] == 17081 && 
b[17082] == 17082 && 
b[17083] == 17083 && 
b[17084] == 17084 && 
b[17085] == 17085 && 
b[17086] == 17086 && 
b[17087] == 17087 && 
b[17088] == 17088 && 
b[17089] == 17089 && 
b[17090] == 17090 && 
b[17091] == 17091 && 
b[17092] == 17092 && 
b[17093] == 17093 && 
b[17094] == 17094 && 
b[17095] == 17095 && 
b[17096] == 17096 && 
b[17097] == 17097 && 
b[17098] == 17098 && 
b[17099] == 17099 && 
b[17100] == 17100 && 
b[17101] == 17101 && 
b[17102] == 17102 && 
b[17103] == 17103 && 
b[17104] == 17104 && 
b[17105] == 17105 && 
b[17106] == 17106 && 
b[17107] == 17107 && 
b[17108] == 17108 && 
b[17109] == 17109 && 
b[17110] == 17110 && 
b[17111] == 17111 && 
b[17112] == 17112 && 
b[17113] == 17113 && 
b[17114] == 17114 && 
b[17115] == 17115 && 
b[17116] == 17116 && 
b[17117] == 17117 && 
b[17118] == 17118 && 
b[17119] == 17119 && 
b[17120] == 17120 && 
b[17121] == 17121 && 
b[17122] == 17122 && 
b[17123] == 17123 && 
b[17124] == 17124 && 
b[17125] == 17125 && 
b[17126] == 17126 && 
b[17127] == 17127 && 
b[17128] == 17128 && 
b[17129] == 17129 && 
b[17130] == 17130 && 
b[17131] == 17131 && 
b[17132] == 17132 && 
b[17133] == 17133 && 
b[17134] == 17134 && 
b[17135] == 17135 && 
b[17136] == 17136 && 
b[17137] == 17137 && 
b[17138] == 17138 && 
b[17139] == 17139 && 
b[17140] == 17140 && 
b[17141] == 17141 && 
b[17142] == 17142 && 
b[17143] == 17143 && 
b[17144] == 17144 && 
b[17145] == 17145 && 
b[17146] == 17146 && 
b[17147] == 17147 && 
b[17148] == 17148 && 
b[17149] == 17149 && 
b[17150] == 17150 && 
b[17151] == 17151 && 
b[17152] == 17152 && 
b[17153] == 17153 && 
b[17154] == 17154 && 
b[17155] == 17155 && 
b[17156] == 17156 && 
b[17157] == 17157 && 
b[17158] == 17158 && 
b[17159] == 17159 && 
b[17160] == 17160 && 
b[17161] == 17161 && 
b[17162] == 17162 && 
b[17163] == 17163 && 
b[17164] == 17164 && 
b[17165] == 17165 && 
b[17166] == 17166 && 
b[17167] == 17167 && 
b[17168] == 17168 && 
b[17169] == 17169 && 
b[17170] == 17170 && 
b[17171] == 17171 && 
b[17172] == 17172 && 
b[17173] == 17173 && 
b[17174] == 17174 && 
b[17175] == 17175 && 
b[17176] == 17176 && 
b[17177] == 17177 && 
b[17178] == 17178 && 
b[17179] == 17179 && 
b[17180] == 17180 && 
b[17181] == 17181 && 
b[17182] == 17182 && 
b[17183] == 17183 && 
b[17184] == 17184 && 
b[17185] == 17185 && 
b[17186] == 17186 && 
b[17187] == 17187 && 
b[17188] == 17188 && 
b[17189] == 17189 && 
b[17190] == 17190 && 
b[17191] == 17191 && 
b[17192] == 17192 && 
b[17193] == 17193 && 
b[17194] == 17194 && 
b[17195] == 17195 && 
b[17196] == 17196 && 
b[17197] == 17197 && 
b[17198] == 17198 && 
b[17199] == 17199 && 
b[17200] == 17200 && 
b[17201] == 17201 && 
b[17202] == 17202 && 
b[17203] == 17203 && 
b[17204] == 17204 && 
b[17205] == 17205 && 
b[17206] == 17206 && 
b[17207] == 17207 && 
b[17208] == 17208 && 
b[17209] == 17209 && 
b[17210] == 17210 && 
b[17211] == 17211 && 
b[17212] == 17212 && 
b[17213] == 17213 && 
b[17214] == 17214 && 
b[17215] == 17215 && 
b[17216] == 17216 && 
b[17217] == 17217 && 
b[17218] == 17218 && 
b[17219] == 17219 && 
b[17220] == 17220 && 
b[17221] == 17221 && 
b[17222] == 17222 && 
b[17223] == 17223 && 
b[17224] == 17224 && 
b[17225] == 17225 && 
b[17226] == 17226 && 
b[17227] == 17227 && 
b[17228] == 17228 && 
b[17229] == 17229 && 
b[17230] == 17230 && 
b[17231] == 17231 && 
b[17232] == 17232 && 
b[17233] == 17233 && 
b[17234] == 17234 && 
b[17235] == 17235 && 
b[17236] == 17236 && 
b[17237] == 17237 && 
b[17238] == 17238 && 
b[17239] == 17239 && 
b[17240] == 17240 && 
b[17241] == 17241 && 
b[17242] == 17242 && 
b[17243] == 17243 && 
b[17244] == 17244 && 
b[17245] == 17245 && 
b[17246] == 17246 && 
b[17247] == 17247 && 
b[17248] == 17248 && 
b[17249] == 17249 && 
b[17250] == 17250 && 
b[17251] == 17251 && 
b[17252] == 17252 && 
b[17253] == 17253 && 
b[17254] == 17254 && 
b[17255] == 17255 && 
b[17256] == 17256 && 
b[17257] == 17257 && 
b[17258] == 17258 && 
b[17259] == 17259 && 
b[17260] == 17260 && 
b[17261] == 17261 && 
b[17262] == 17262 && 
b[17263] == 17263 && 
b[17264] == 17264 && 
b[17265] == 17265 && 
b[17266] == 17266 && 
b[17267] == 17267 && 
b[17268] == 17268 && 
b[17269] == 17269 && 
b[17270] == 17270 && 
b[17271] == 17271 && 
b[17272] == 17272 && 
b[17273] == 17273 && 
b[17274] == 17274 && 
b[17275] == 17275 && 
b[17276] == 17276 && 
b[17277] == 17277 && 
b[17278] == 17278 && 
b[17279] == 17279 && 
b[17280] == 17280 && 
b[17281] == 17281 && 
b[17282] == 17282 && 
b[17283] == 17283 && 
b[17284] == 17284 && 
b[17285] == 17285 && 
b[17286] == 17286 && 
b[17287] == 17287 && 
b[17288] == 17288 && 
b[17289] == 17289 && 
b[17290] == 17290 && 
b[17291] == 17291 && 
b[17292] == 17292 && 
b[17293] == 17293 && 
b[17294] == 17294 && 
b[17295] == 17295 && 
b[17296] == 17296 && 
b[17297] == 17297 && 
b[17298] == 17298 && 
b[17299] == 17299 && 
b[17300] == 17300 && 
b[17301] == 17301 && 
b[17302] == 17302 && 
b[17303] == 17303 && 
b[17304] == 17304 && 
b[17305] == 17305 && 
b[17306] == 17306 && 
b[17307] == 17307 && 
b[17308] == 17308 && 
b[17309] == 17309 && 
b[17310] == 17310 && 
b[17311] == 17311 && 
b[17312] == 17312 && 
b[17313] == 17313 && 
b[17314] == 17314 && 
b[17315] == 17315 && 
b[17316] == 17316 && 
b[17317] == 17317 && 
b[17318] == 17318 && 
b[17319] == 17319 && 
b[17320] == 17320 && 
b[17321] == 17321 && 
b[17322] == 17322 && 
b[17323] == 17323 && 
b[17324] == 17324 && 
b[17325] == 17325 && 
b[17326] == 17326 && 
b[17327] == 17327 && 
b[17328] == 17328 && 
b[17329] == 17329 && 
b[17330] == 17330 && 
b[17331] == 17331 && 
b[17332] == 17332 && 
b[17333] == 17333 && 
b[17334] == 17334 && 
b[17335] == 17335 && 
b[17336] == 17336 && 
b[17337] == 17337 && 
b[17338] == 17338 && 
b[17339] == 17339 && 
b[17340] == 17340 && 
b[17341] == 17341 && 
b[17342] == 17342 && 
b[17343] == 17343 && 
b[17344] == 17344 && 
b[17345] == 17345 && 
b[17346] == 17346 && 
b[17347] == 17347 && 
b[17348] == 17348 && 
b[17349] == 17349 && 
b[17350] == 17350 && 
b[17351] == 17351 && 
b[17352] == 17352 && 
b[17353] == 17353 && 
b[17354] == 17354 && 
b[17355] == 17355 && 
b[17356] == 17356 && 
b[17357] == 17357 && 
b[17358] == 17358 && 
b[17359] == 17359 && 
b[17360] == 17360 && 
b[17361] == 17361 && 
b[17362] == 17362 && 
b[17363] == 17363 && 
b[17364] == 17364 && 
b[17365] == 17365 && 
b[17366] == 17366 && 
b[17367] == 17367 && 
b[17368] == 17368 && 
b[17369] == 17369 && 
b[17370] == 17370 && 
b[17371] == 17371 && 
b[17372] == 17372 && 
b[17373] == 17373 && 
b[17374] == 17374 && 
b[17375] == 17375 && 
b[17376] == 17376 && 
b[17377] == 17377 && 
b[17378] == 17378 && 
b[17379] == 17379 && 
b[17380] == 17380 && 
b[17381] == 17381 && 
b[17382] == 17382 && 
b[17383] == 17383 && 
b[17384] == 17384 && 
b[17385] == 17385 && 
b[17386] == 17386 && 
b[17387] == 17387 && 
b[17388] == 17388 && 
b[17389] == 17389 && 
b[17390] == 17390 && 
b[17391] == 17391 && 
b[17392] == 17392 && 
b[17393] == 17393 && 
b[17394] == 17394 && 
b[17395] == 17395 && 
b[17396] == 17396 && 
b[17397] == 17397 && 
b[17398] == 17398 && 
b[17399] == 17399 && 
b[17400] == 17400 && 
b[17401] == 17401 && 
b[17402] == 17402 && 
b[17403] == 17403 && 
b[17404] == 17404 && 
b[17405] == 17405 && 
b[17406] == 17406 && 
b[17407] == 17407 && 
b[17408] == 17408 && 
b[17409] == 17409 && 
b[17410] == 17410 && 
b[17411] == 17411 && 
b[17412] == 17412 && 
b[17413] == 17413 && 
b[17414] == 17414 && 
b[17415] == 17415 && 
b[17416] == 17416 && 
b[17417] == 17417 && 
b[17418] == 17418 && 
b[17419] == 17419 && 
b[17420] == 17420 && 
b[17421] == 17421 && 
b[17422] == 17422 && 
b[17423] == 17423 && 
b[17424] == 17424 && 
b[17425] == 17425 && 
b[17426] == 17426 && 
b[17427] == 17427 && 
b[17428] == 17428 && 
b[17429] == 17429 && 
b[17430] == 17430 && 
b[17431] == 17431 && 
b[17432] == 17432 && 
b[17433] == 17433 && 
b[17434] == 17434 && 
b[17435] == 17435 && 
b[17436] == 17436 && 
b[17437] == 17437 && 
b[17438] == 17438 && 
b[17439] == 17439 && 
b[17440] == 17440 && 
b[17441] == 17441 && 
b[17442] == 17442 && 
b[17443] == 17443 && 
b[17444] == 17444 && 
b[17445] == 17445 && 
b[17446] == 17446 && 
b[17447] == 17447 && 
b[17448] == 17448 && 
b[17449] == 17449 && 
b[17450] == 17450 && 
b[17451] == 17451 && 
b[17452] == 17452 && 
b[17453] == 17453 && 
b[17454] == 17454 && 
b[17455] == 17455 && 
b[17456] == 17456 && 
b[17457] == 17457 && 
b[17458] == 17458 && 
b[17459] == 17459 && 
b[17460] == 17460 && 
b[17461] == 17461 && 
b[17462] == 17462 && 
b[17463] == 17463 && 
b[17464] == 17464 && 
b[17465] == 17465 && 
b[17466] == 17466 && 
b[17467] == 17467 && 
b[17468] == 17468 && 
b[17469] == 17469 && 
b[17470] == 17470 && 
b[17471] == 17471 && 
b[17472] == 17472 && 
b[17473] == 17473 && 
b[17474] == 17474 && 
b[17475] == 17475 && 
b[17476] == 17476 && 
b[17477] == 17477 && 
b[17478] == 17478 && 
b[17479] == 17479 && 
b[17480] == 17480 && 
b[17481] == 17481 && 
b[17482] == 17482 && 
b[17483] == 17483 && 
b[17484] == 17484 && 
b[17485] == 17485 && 
b[17486] == 17486 && 
b[17487] == 17487 && 
b[17488] == 17488 && 
b[17489] == 17489 && 
b[17490] == 17490 && 
b[17491] == 17491 && 
b[17492] == 17492 && 
b[17493] == 17493 && 
b[17494] == 17494 && 
b[17495] == 17495 && 
b[17496] == 17496 && 
b[17497] == 17497 && 
b[17498] == 17498 && 
b[17499] == 17499 && 
b[17500] == 17500 && 
b[17501] == 17501 && 
b[17502] == 17502 && 
b[17503] == 17503 && 
b[17504] == 17504 && 
b[17505] == 17505 && 
b[17506] == 17506 && 
b[17507] == 17507 && 
b[17508] == 17508 && 
b[17509] == 17509 && 
b[17510] == 17510 && 
b[17511] == 17511 && 
b[17512] == 17512 && 
b[17513] == 17513 && 
b[17514] == 17514 && 
b[17515] == 17515 && 
b[17516] == 17516 && 
b[17517] == 17517 && 
b[17518] == 17518 && 
b[17519] == 17519 && 
b[17520] == 17520 && 
b[17521] == 17521 && 
b[17522] == 17522 && 
b[17523] == 17523 && 
b[17524] == 17524 && 
b[17525] == 17525 && 
b[17526] == 17526 && 
b[17527] == 17527 && 
b[17528] == 17528 && 
b[17529] == 17529 && 
b[17530] == 17530 && 
b[17531] == 17531 && 
b[17532] == 17532 && 
b[17533] == 17533 && 
b[17534] == 17534 && 
b[17535] == 17535 && 
b[17536] == 17536 && 
b[17537] == 17537 && 
b[17538] == 17538 && 
b[17539] == 17539 && 
b[17540] == 17540 && 
b[17541] == 17541 && 
b[17542] == 17542 && 
b[17543] == 17543 && 
b[17544] == 17544 && 
b[17545] == 17545 && 
b[17546] == 17546 && 
b[17547] == 17547 && 
b[17548] == 17548 && 
b[17549] == 17549 && 
b[17550] == 17550 && 
b[17551] == 17551 && 
b[17552] == 17552 && 
b[17553] == 17553 && 
b[17554] == 17554 && 
b[17555] == 17555 && 
b[17556] == 17556 && 
b[17557] == 17557 && 
b[17558] == 17558 && 
b[17559] == 17559 && 
b[17560] == 17560 && 
b[17561] == 17561 && 
b[17562] == 17562 && 
b[17563] == 17563 && 
b[17564] == 17564 && 
b[17565] == 17565 && 
b[17566] == 17566 && 
b[17567] == 17567 && 
b[17568] == 17568 && 
b[17569] == 17569 && 
b[17570] == 17570 && 
b[17571] == 17571 && 
b[17572] == 17572 && 
b[17573] == 17573 && 
b[17574] == 17574 && 
b[17575] == 17575 && 
b[17576] == 17576 && 
b[17577] == 17577 && 
b[17578] == 17578 && 
b[17579] == 17579 && 
b[17580] == 17580 && 
b[17581] == 17581 && 
b[17582] == 17582 && 
b[17583] == 17583 && 
b[17584] == 17584 && 
b[17585] == 17585 && 
b[17586] == 17586 && 
b[17587] == 17587 && 
b[17588] == 17588 && 
b[17589] == 17589 && 
b[17590] == 17590 && 
b[17591] == 17591 && 
b[17592] == 17592 && 
b[17593] == 17593 && 
b[17594] == 17594 && 
b[17595] == 17595 && 
b[17596] == 17596 && 
b[17597] == 17597 && 
b[17598] == 17598 && 
b[17599] == 17599 && 
b[17600] == 17600 && 
b[17601] == 17601 && 
b[17602] == 17602 && 
b[17603] == 17603 && 
b[17604] == 17604 && 
b[17605] == 17605 && 
b[17606] == 17606 && 
b[17607] == 17607 && 
b[17608] == 17608 && 
b[17609] == 17609 && 
b[17610] == 17610 && 
b[17611] == 17611 && 
b[17612] == 17612 && 
b[17613] == 17613 && 
b[17614] == 17614 && 
b[17615] == 17615 && 
b[17616] == 17616 && 
b[17617] == 17617 && 
b[17618] == 17618 && 
b[17619] == 17619 && 
b[17620] == 17620 && 
b[17621] == 17621 && 
b[17622] == 17622 && 
b[17623] == 17623 && 
b[17624] == 17624 && 
b[17625] == 17625 && 
b[17626] == 17626 && 
b[17627] == 17627 && 
b[17628] == 17628 && 
b[17629] == 17629 && 
b[17630] == 17630 && 
b[17631] == 17631 && 
b[17632] == 17632 && 
b[17633] == 17633 && 
b[17634] == 17634 && 
b[17635] == 17635 && 
b[17636] == 17636 && 
b[17637] == 17637 && 
b[17638] == 17638 && 
b[17639] == 17639 && 
b[17640] == 17640 && 
b[17641] == 17641 && 
b[17642] == 17642 && 
b[17643] == 17643 && 
b[17644] == 17644 && 
b[17645] == 17645 && 
b[17646] == 17646 && 
b[17647] == 17647 && 
b[17648] == 17648 && 
b[17649] == 17649 && 
b[17650] == 17650 && 
b[17651] == 17651 && 
b[17652] == 17652 && 
b[17653] == 17653 && 
b[17654] == 17654 && 
b[17655] == 17655 && 
b[17656] == 17656 && 
b[17657] == 17657 && 
b[17658] == 17658 && 
b[17659] == 17659 && 
b[17660] == 17660 && 
b[17661] == 17661 && 
b[17662] == 17662 && 
b[17663] == 17663 && 
b[17664] == 17664 && 
b[17665] == 17665 && 
b[17666] == 17666 && 
b[17667] == 17667 && 
b[17668] == 17668 && 
b[17669] == 17669 && 
b[17670] == 17670 && 
b[17671] == 17671 && 
b[17672] == 17672 && 
b[17673] == 17673 && 
b[17674] == 17674 && 
b[17675] == 17675 && 
b[17676] == 17676 && 
b[17677] == 17677 && 
b[17678] == 17678 && 
b[17679] == 17679 && 
b[17680] == 17680 && 
b[17681] == 17681 && 
b[17682] == 17682 && 
b[17683] == 17683 && 
b[17684] == 17684 && 
b[17685] == 17685 && 
b[17686] == 17686 && 
b[17687] == 17687 && 
b[17688] == 17688 && 
b[17689] == 17689 && 
b[17690] == 17690 && 
b[17691] == 17691 && 
b[17692] == 17692 && 
b[17693] == 17693 && 
b[17694] == 17694 && 
b[17695] == 17695 && 
b[17696] == 17696 && 
b[17697] == 17697 && 
b[17698] == 17698 && 
b[17699] == 17699 && 
b[17700] == 17700 && 
b[17701] == 17701 && 
b[17702] == 17702 && 
b[17703] == 17703 && 
b[17704] == 17704 && 
b[17705] == 17705 && 
b[17706] == 17706 && 
b[17707] == 17707 && 
b[17708] == 17708 && 
b[17709] == 17709 && 
b[17710] == 17710 && 
b[17711] == 17711 && 
b[17712] == 17712 && 
b[17713] == 17713 && 
b[17714] == 17714 && 
b[17715] == 17715 && 
b[17716] == 17716 && 
b[17717] == 17717 && 
b[17718] == 17718 && 
b[17719] == 17719 && 
b[17720] == 17720 && 
b[17721] == 17721 && 
b[17722] == 17722 && 
b[17723] == 17723 && 
b[17724] == 17724 && 
b[17725] == 17725 && 
b[17726] == 17726 && 
b[17727] == 17727 && 
b[17728] == 17728 && 
b[17729] == 17729 && 
b[17730] == 17730 && 
b[17731] == 17731 && 
b[17732] == 17732 && 
b[17733] == 17733 && 
b[17734] == 17734 && 
b[17735] == 17735 && 
b[17736] == 17736 && 
b[17737] == 17737 && 
b[17738] == 17738 && 
b[17739] == 17739 && 
b[17740] == 17740 && 
b[17741] == 17741 && 
b[17742] == 17742 && 
b[17743] == 17743 && 
b[17744] == 17744 && 
b[17745] == 17745 && 
b[17746] == 17746 && 
b[17747] == 17747 && 
b[17748] == 17748 && 
b[17749] == 17749 && 
b[17750] == 17750 && 
b[17751] == 17751 && 
b[17752] == 17752 && 
b[17753] == 17753 && 
b[17754] == 17754 && 
b[17755] == 17755 && 
b[17756] == 17756 && 
b[17757] == 17757 && 
b[17758] == 17758 && 
b[17759] == 17759 && 
b[17760] == 17760 && 
b[17761] == 17761 && 
b[17762] == 17762 && 
b[17763] == 17763 && 
b[17764] == 17764 && 
b[17765] == 17765 && 
b[17766] == 17766 && 
b[17767] == 17767 && 
b[17768] == 17768 && 
b[17769] == 17769 && 
b[17770] == 17770 && 
b[17771] == 17771 && 
b[17772] == 17772 && 
b[17773] == 17773 && 
b[17774] == 17774 && 
b[17775] == 17775 && 
b[17776] == 17776 && 
b[17777] == 17777 && 
b[17778] == 17778 && 
b[17779] == 17779 && 
b[17780] == 17780 && 
b[17781] == 17781 && 
b[17782] == 17782 && 
b[17783] == 17783 && 
b[17784] == 17784 && 
b[17785] == 17785 && 
b[17786] == 17786 && 
b[17787] == 17787 && 
b[17788] == 17788 && 
b[17789] == 17789 && 
b[17790] == 17790 && 
b[17791] == 17791 && 
b[17792] == 17792 && 
b[17793] == 17793 && 
b[17794] == 17794 && 
b[17795] == 17795 && 
b[17796] == 17796 && 
b[17797] == 17797 && 
b[17798] == 17798 && 
b[17799] == 17799 && 
b[17800] == 17800 && 
b[17801] == 17801 && 
b[17802] == 17802 && 
b[17803] == 17803 && 
b[17804] == 17804 && 
b[17805] == 17805 && 
b[17806] == 17806 && 
b[17807] == 17807 && 
b[17808] == 17808 && 
b[17809] == 17809 && 
b[17810] == 17810 && 
b[17811] == 17811 && 
b[17812] == 17812 && 
b[17813] == 17813 && 
b[17814] == 17814 && 
b[17815] == 17815 && 
b[17816] == 17816 && 
b[17817] == 17817 && 
b[17818] == 17818 && 
b[17819] == 17819 && 
b[17820] == 17820 && 
b[17821] == 17821 && 
b[17822] == 17822 && 
b[17823] == 17823 && 
b[17824] == 17824 && 
b[17825] == 17825 && 
b[17826] == 17826 && 
b[17827] == 17827 && 
b[17828] == 17828 && 
b[17829] == 17829 && 
b[17830] == 17830 && 
b[17831] == 17831 && 
b[17832] == 17832 && 
b[17833] == 17833 && 
b[17834] == 17834 && 
b[17835] == 17835 && 
b[17836] == 17836 && 
b[17837] == 17837 && 
b[17838] == 17838 && 
b[17839] == 17839 && 
b[17840] == 17840 && 
b[17841] == 17841 && 
b[17842] == 17842 && 
b[17843] == 17843 && 
b[17844] == 17844 && 
b[17845] == 17845 && 
b[17846] == 17846 && 
b[17847] == 17847 && 
b[17848] == 17848 && 
b[17849] == 17849 && 
b[17850] == 17850 && 
b[17851] == 17851 && 
b[17852] == 17852 && 
b[17853] == 17853 && 
b[17854] == 17854 && 
b[17855] == 17855 && 
b[17856] == 17856 && 
b[17857] == 17857 && 
b[17858] == 17858 && 
b[17859] == 17859 && 
b[17860] == 17860 && 
b[17861] == 17861 && 
b[17862] == 17862 && 
b[17863] == 17863 && 
b[17864] == 17864 && 
b[17865] == 17865 && 
b[17866] == 17866 && 
b[17867] == 17867 && 
b[17868] == 17868 && 
b[17869] == 17869 && 
b[17870] == 17870 && 
b[17871] == 17871 && 
b[17872] == 17872 && 
b[17873] == 17873 && 
b[17874] == 17874 && 
b[17875] == 17875 && 
b[17876] == 17876 && 
b[17877] == 17877 && 
b[17878] == 17878 && 
b[17879] == 17879 && 
b[17880] == 17880 && 
b[17881] == 17881 && 
b[17882] == 17882 && 
b[17883] == 17883 && 
b[17884] == 17884 && 
b[17885] == 17885 && 
b[17886] == 17886 && 
b[17887] == 17887 && 
b[17888] == 17888 && 
b[17889] == 17889 && 
b[17890] == 17890 && 
b[17891] == 17891 && 
b[17892] == 17892 && 
b[17893] == 17893 && 
b[17894] == 17894 && 
b[17895] == 17895 && 
b[17896] == 17896 && 
b[17897] == 17897 && 
b[17898] == 17898 && 
b[17899] == 17899 && 
b[17900] == 17900 && 
b[17901] == 17901 && 
b[17902] == 17902 && 
b[17903] == 17903 && 
b[17904] == 17904 && 
b[17905] == 17905 && 
b[17906] == 17906 && 
b[17907] == 17907 && 
b[17908] == 17908 && 
b[17909] == 17909 && 
b[17910] == 17910 && 
b[17911] == 17911 && 
b[17912] == 17912 && 
b[17913] == 17913 && 
b[17914] == 17914 && 
b[17915] == 17915 && 
b[17916] == 17916 && 
b[17917] == 17917 && 
b[17918] == 17918 && 
b[17919] == 17919 && 
b[17920] == 17920 && 
b[17921] == 17921 && 
b[17922] == 17922 && 
b[17923] == 17923 && 
b[17924] == 17924 && 
b[17925] == 17925 && 
b[17926] == 17926 && 
b[17927] == 17927 && 
b[17928] == 17928 && 
b[17929] == 17929 && 
b[17930] == 17930 && 
b[17931] == 17931 && 
b[17932] == 17932 && 
b[17933] == 17933 && 
b[17934] == 17934 && 
b[17935] == 17935 && 
b[17936] == 17936 && 
b[17937] == 17937 && 
b[17938] == 17938 && 
b[17939] == 17939 && 
b[17940] == 17940 && 
b[17941] == 17941 && 
b[17942] == 17942 && 
b[17943] == 17943 && 
b[17944] == 17944 && 
b[17945] == 17945 && 
b[17946] == 17946 && 
b[17947] == 17947 && 
b[17948] == 17948 && 
b[17949] == 17949 && 
b[17950] == 17950 && 
b[17951] == 17951 && 
b[17952] == 17952 && 
b[17953] == 17953 && 
b[17954] == 17954 && 
b[17955] == 17955 && 
b[17956] == 17956 && 
b[17957] == 17957 && 
b[17958] == 17958 && 
b[17959] == 17959 && 
b[17960] == 17960 && 
b[17961] == 17961 && 
b[17962] == 17962 && 
b[17963] == 17963 && 
b[17964] == 17964 && 
b[17965] == 17965 && 
b[17966] == 17966 && 
b[17967] == 17967 && 
b[17968] == 17968 && 
b[17969] == 17969 && 
b[17970] == 17970 && 
b[17971] == 17971 && 
b[17972] == 17972 && 
b[17973] == 17973 && 
b[17974] == 17974 && 
b[17975] == 17975 && 
b[17976] == 17976 && 
b[17977] == 17977 && 
b[17978] == 17978 && 
b[17979] == 17979 && 
b[17980] == 17980 && 
b[17981] == 17981 && 
b[17982] == 17982 && 
b[17983] == 17983 && 
b[17984] == 17984 && 
b[17985] == 17985 && 
b[17986] == 17986 && 
b[17987] == 17987 && 
b[17988] == 17988 && 
b[17989] == 17989 && 
b[17990] == 17990 && 
b[17991] == 17991 && 
b[17992] == 17992 && 
b[17993] == 17993 && 
b[17994] == 17994 && 
b[17995] == 17995 && 
b[17996] == 17996 && 
b[17997] == 17997 && 
b[17998] == 17998 && 
b[17999] == 17999 && 
b[18000] == 18000 && 
b[18001] == 18001 && 
b[18002] == 18002 && 
b[18003] == 18003 && 
b[18004] == 18004 && 
b[18005] == 18005 && 
b[18006] == 18006 && 
b[18007] == 18007 && 
b[18008] == 18008 && 
b[18009] == 18009 && 
b[18010] == 18010 && 
b[18011] == 18011 && 
b[18012] == 18012 && 
b[18013] == 18013 && 
b[18014] == 18014 && 
b[18015] == 18015 && 
b[18016] == 18016 && 
b[18017] == 18017 && 
b[18018] == 18018 && 
b[18019] == 18019 && 
b[18020] == 18020 && 
b[18021] == 18021 && 
b[18022] == 18022 && 
b[18023] == 18023 && 
b[18024] == 18024 && 
b[18025] == 18025 && 
b[18026] == 18026 && 
b[18027] == 18027 && 
b[18028] == 18028 && 
b[18029] == 18029 && 
b[18030] == 18030 && 
b[18031] == 18031 && 
b[18032] == 18032 && 
b[18033] == 18033 && 
b[18034] == 18034 && 
b[18035] == 18035 && 
b[18036] == 18036 && 
b[18037] == 18037 && 
b[18038] == 18038 && 
b[18039] == 18039 && 
b[18040] == 18040 && 
b[18041] == 18041 && 
b[18042] == 18042 && 
b[18043] == 18043 && 
b[18044] == 18044 && 
b[18045] == 18045 && 
b[18046] == 18046 && 
b[18047] == 18047 && 
b[18048] == 18048 && 
b[18049] == 18049 && 
b[18050] == 18050 && 
b[18051] == 18051 && 
b[18052] == 18052 && 
b[18053] == 18053 && 
b[18054] == 18054 && 
b[18055] == 18055 && 
b[18056] == 18056 && 
b[18057] == 18057 && 
b[18058] == 18058 && 
b[18059] == 18059 && 
b[18060] == 18060 && 
b[18061] == 18061 && 
b[18062] == 18062 && 
b[18063] == 18063 && 
b[18064] == 18064 && 
b[18065] == 18065 && 
b[18066] == 18066 && 
b[18067] == 18067 && 
b[18068] == 18068 && 
b[18069] == 18069 && 
b[18070] == 18070 && 
b[18071] == 18071 && 
b[18072] == 18072 && 
b[18073] == 18073 && 
b[18074] == 18074 && 
b[18075] == 18075 && 
b[18076] == 18076 && 
b[18077] == 18077 && 
b[18078] == 18078 && 
b[18079] == 18079 && 
b[18080] == 18080 && 
b[18081] == 18081 && 
b[18082] == 18082 && 
b[18083] == 18083 && 
b[18084] == 18084 && 
b[18085] == 18085 && 
b[18086] == 18086 && 
b[18087] == 18087 && 
b[18088] == 18088 && 
b[18089] == 18089 && 
b[18090] == 18090 && 
b[18091] == 18091 && 
b[18092] == 18092 && 
b[18093] == 18093 && 
b[18094] == 18094 && 
b[18095] == 18095 && 
b[18096] == 18096 && 
b[18097] == 18097 && 
b[18098] == 18098 && 
b[18099] == 18099 && 
b[18100] == 18100 && 
b[18101] == 18101 && 
b[18102] == 18102 && 
b[18103] == 18103 && 
b[18104] == 18104 && 
b[18105] == 18105 && 
b[18106] == 18106 && 
b[18107] == 18107 && 
b[18108] == 18108 && 
b[18109] == 18109 && 
b[18110] == 18110 && 
b[18111] == 18111 && 
b[18112] == 18112 && 
b[18113] == 18113 && 
b[18114] == 18114 && 
b[18115] == 18115 && 
b[18116] == 18116 && 
b[18117] == 18117 && 
b[18118] == 18118 && 
b[18119] == 18119 && 
b[18120] == 18120 && 
b[18121] == 18121 && 
b[18122] == 18122 && 
b[18123] == 18123 && 
b[18124] == 18124 && 
b[18125] == 18125 && 
b[18126] == 18126 && 
b[18127] == 18127 && 
b[18128] == 18128 && 
b[18129] == 18129 && 
b[18130] == 18130 && 
b[18131] == 18131 && 
b[18132] == 18132 && 
b[18133] == 18133 && 
b[18134] == 18134 && 
b[18135] == 18135 && 
b[18136] == 18136 && 
b[18137] == 18137 && 
b[18138] == 18138 && 
b[18139] == 18139 && 
b[18140] == 18140 && 
b[18141] == 18141 && 
b[18142] == 18142 && 
b[18143] == 18143 && 
b[18144] == 18144 && 
b[18145] == 18145 && 
b[18146] == 18146 && 
b[18147] == 18147 && 
b[18148] == 18148 && 
b[18149] == 18149 && 
b[18150] == 18150 && 
b[18151] == 18151 && 
b[18152] == 18152 && 
b[18153] == 18153 && 
b[18154] == 18154 && 
b[18155] == 18155 && 
b[18156] == 18156 && 
b[18157] == 18157 && 
b[18158] == 18158 && 
b[18159] == 18159 && 
b[18160] == 18160 && 
b[18161] == 18161 && 
b[18162] == 18162 && 
b[18163] == 18163 && 
b[18164] == 18164 && 
b[18165] == 18165 && 
b[18166] == 18166 && 
b[18167] == 18167 && 
b[18168] == 18168 && 
b[18169] == 18169 && 
b[18170] == 18170 && 
b[18171] == 18171 && 
b[18172] == 18172 && 
b[18173] == 18173 && 
b[18174] == 18174 && 
b[18175] == 18175 && 
b[18176] == 18176 && 
b[18177] == 18177 && 
b[18178] == 18178 && 
b[18179] == 18179 && 
b[18180] == 18180 && 
b[18181] == 18181 && 
b[18182] == 18182 && 
b[18183] == 18183 && 
b[18184] == 18184 && 
b[18185] == 18185 && 
b[18186] == 18186 && 
b[18187] == 18187 && 
b[18188] == 18188 && 
b[18189] == 18189 && 
b[18190] == 18190 && 
b[18191] == 18191 && 
b[18192] == 18192 && 
b[18193] == 18193 && 
b[18194] == 18194 && 
b[18195] == 18195 && 
b[18196] == 18196 && 
b[18197] == 18197 && 
b[18198] == 18198 && 
b[18199] == 18199 && 
b[18200] == 18200 && 
b[18201] == 18201 && 
b[18202] == 18202 && 
b[18203] == 18203 && 
b[18204] == 18204 && 
b[18205] == 18205 && 
b[18206] == 18206 && 
b[18207] == 18207 && 
b[18208] == 18208 && 
b[18209] == 18209 && 
b[18210] == 18210 && 
b[18211] == 18211 && 
b[18212] == 18212 && 
b[18213] == 18213 && 
b[18214] == 18214 && 
b[18215] == 18215 && 
b[18216] == 18216 && 
b[18217] == 18217 && 
b[18218] == 18218 && 
b[18219] == 18219 && 
b[18220] == 18220 && 
b[18221] == 18221 && 
b[18222] == 18222 && 
b[18223] == 18223 && 
b[18224] == 18224 && 
b[18225] == 18225 && 
b[18226] == 18226 && 
b[18227] == 18227 && 
b[18228] == 18228 && 
b[18229] == 18229 && 
b[18230] == 18230 && 
b[18231] == 18231 && 
b[18232] == 18232 && 
b[18233] == 18233 && 
b[18234] == 18234 && 
b[18235] == 18235 && 
b[18236] == 18236 && 
b[18237] == 18237 && 
b[18238] == 18238 && 
b[18239] == 18239 && 
b[18240] == 18240 && 
b[18241] == 18241 && 
b[18242] == 18242 && 
b[18243] == 18243 && 
b[18244] == 18244 && 
b[18245] == 18245 && 
b[18246] == 18246 && 
b[18247] == 18247 && 
b[18248] == 18248 && 
b[18249] == 18249 && 
b[18250] == 18250 && 
b[18251] == 18251 && 
b[18252] == 18252 && 
b[18253] == 18253 && 
b[18254] == 18254 && 
b[18255] == 18255 && 
b[18256] == 18256 && 
b[18257] == 18257 && 
b[18258] == 18258 && 
b[18259] == 18259 && 
b[18260] == 18260 && 
b[18261] == 18261 && 
b[18262] == 18262 && 
b[18263] == 18263 && 
b[18264] == 18264 && 
b[18265] == 18265 && 
b[18266] == 18266 && 
b[18267] == 18267 && 
b[18268] == 18268 && 
b[18269] == 18269 && 
b[18270] == 18270 && 
b[18271] == 18271 && 
b[18272] == 18272 && 
b[18273] == 18273 && 
b[18274] == 18274 && 
b[18275] == 18275 && 
b[18276] == 18276 && 
b[18277] == 18277 && 
b[18278] == 18278 && 
b[18279] == 18279 && 
b[18280] == 18280 && 
b[18281] == 18281 && 
b[18282] == 18282 && 
b[18283] == 18283 && 
b[18284] == 18284 && 
b[18285] == 18285 && 
b[18286] == 18286 && 
b[18287] == 18287 && 
b[18288] == 18288 && 
b[18289] == 18289 && 
b[18290] == 18290 && 
b[18291] == 18291 && 
b[18292] == 18292 && 
b[18293] == 18293 && 
b[18294] == 18294 && 
b[18295] == 18295 && 
b[18296] == 18296 && 
b[18297] == 18297 && 
b[18298] == 18298 && 
b[18299] == 18299 && 
b[18300] == 18300 && 
b[18301] == 18301 && 
b[18302] == 18302 && 
b[18303] == 18303 && 
b[18304] == 18304 && 
b[18305] == 18305 && 
b[18306] == 18306 && 
b[18307] == 18307 && 
b[18308] == 18308 && 
b[18309] == 18309 && 
b[18310] == 18310 && 
b[18311] == 18311 && 
b[18312] == 18312 && 
b[18313] == 18313 && 
b[18314] == 18314 && 
b[18315] == 18315 && 
b[18316] == 18316 && 
b[18317] == 18317 && 
b[18318] == 18318 && 
b[18319] == 18319 && 
b[18320] == 18320 && 
b[18321] == 18321 && 
b[18322] == 18322 && 
b[18323] == 18323 && 
b[18324] == 18324 && 
b[18325] == 18325 && 
b[18326] == 18326 && 
b[18327] == 18327 && 
b[18328] == 18328 && 
b[18329] == 18329 && 
b[18330] == 18330 && 
b[18331] == 18331 && 
b[18332] == 18332 && 
b[18333] == 18333 && 
b[18334] == 18334 && 
b[18335] == 18335 && 
b[18336] == 18336 && 
b[18337] == 18337 && 
b[18338] == 18338 && 
b[18339] == 18339 && 
b[18340] == 18340 && 
b[18341] == 18341 && 
b[18342] == 18342 && 
b[18343] == 18343 && 
b[18344] == 18344 && 
b[18345] == 18345 && 
b[18346] == 18346 && 
b[18347] == 18347 && 
b[18348] == 18348 && 
b[18349] == 18349 && 
b[18350] == 18350 && 
b[18351] == 18351 && 
b[18352] == 18352 && 
b[18353] == 18353 && 
b[18354] == 18354 && 
b[18355] == 18355 && 
b[18356] == 18356 && 
b[18357] == 18357 && 
b[18358] == 18358 && 
b[18359] == 18359 && 
b[18360] == 18360 && 
b[18361] == 18361 && 
b[18362] == 18362 && 
b[18363] == 18363 && 
b[18364] == 18364 && 
b[18365] == 18365 && 
b[18366] == 18366 && 
b[18367] == 18367 && 
b[18368] == 18368 && 
b[18369] == 18369 && 
b[18370] == 18370 && 
b[18371] == 18371 && 
b[18372] == 18372 && 
b[18373] == 18373 && 
b[18374] == 18374 && 
b[18375] == 18375 && 
b[18376] == 18376 && 
b[18377] == 18377 && 
b[18378] == 18378 && 
b[18379] == 18379 && 
b[18380] == 18380 && 
b[18381] == 18381 && 
b[18382] == 18382 && 
b[18383] == 18383 && 
b[18384] == 18384 && 
b[18385] == 18385 && 
b[18386] == 18386 && 
b[18387] == 18387 && 
b[18388] == 18388 && 
b[18389] == 18389 && 
b[18390] == 18390 && 
b[18391] == 18391 && 
b[18392] == 18392 && 
b[18393] == 18393 && 
b[18394] == 18394 && 
b[18395] == 18395 && 
b[18396] == 18396 && 
b[18397] == 18397 && 
b[18398] == 18398 && 
b[18399] == 18399 && 
b[18400] == 18400 && 
b[18401] == 18401 && 
b[18402] == 18402 && 
b[18403] == 18403 && 
b[18404] == 18404 && 
b[18405] == 18405 && 
b[18406] == 18406 && 
b[18407] == 18407 && 
b[18408] == 18408 && 
b[18409] == 18409 && 
b[18410] == 18410 && 
b[18411] == 18411 && 
b[18412] == 18412 && 
b[18413] == 18413 && 
b[18414] == 18414 && 
b[18415] == 18415 && 
b[18416] == 18416 && 
b[18417] == 18417 && 
b[18418] == 18418 && 
b[18419] == 18419 && 
b[18420] == 18420 && 
b[18421] == 18421 && 
b[18422] == 18422 && 
b[18423] == 18423 && 
b[18424] == 18424 && 
b[18425] == 18425 && 
b[18426] == 18426 && 
b[18427] == 18427 && 
b[18428] == 18428 && 
b[18429] == 18429 && 
b[18430] == 18430 && 
b[18431] == 18431 && 
b[18432] == 18432 && 
b[18433] == 18433 && 
b[18434] == 18434 && 
b[18435] == 18435 && 
b[18436] == 18436 && 
b[18437] == 18437 && 
b[18438] == 18438 && 
b[18439] == 18439 && 
b[18440] == 18440 && 
b[18441] == 18441 && 
b[18442] == 18442 && 
b[18443] == 18443 && 
b[18444] == 18444 && 
b[18445] == 18445 && 
b[18446] == 18446 && 
b[18447] == 18447 && 
b[18448] == 18448 && 
b[18449] == 18449 && 
b[18450] == 18450 && 
b[18451] == 18451 && 
b[18452] == 18452 && 
b[18453] == 18453 && 
b[18454] == 18454 && 
b[18455] == 18455 && 
b[18456] == 18456 && 
b[18457] == 18457 && 
b[18458] == 18458 && 
b[18459] == 18459 && 
b[18460] == 18460 && 
b[18461] == 18461 && 
b[18462] == 18462 && 
b[18463] == 18463 && 
b[18464] == 18464 && 
b[18465] == 18465 && 
b[18466] == 18466 && 
b[18467] == 18467 && 
b[18468] == 18468 && 
b[18469] == 18469 && 
b[18470] == 18470 && 
b[18471] == 18471 && 
b[18472] == 18472 && 
b[18473] == 18473 && 
b[18474] == 18474 && 
b[18475] == 18475 && 
b[18476] == 18476 && 
b[18477] == 18477 && 
b[18478] == 18478 && 
b[18479] == 18479 && 
b[18480] == 18480 && 
b[18481] == 18481 && 
b[18482] == 18482 && 
b[18483] == 18483 && 
b[18484] == 18484 && 
b[18485] == 18485 && 
b[18486] == 18486 && 
b[18487] == 18487 && 
b[18488] == 18488 && 
b[18489] == 18489 && 
b[18490] == 18490 && 
b[18491] == 18491 && 
b[18492] == 18492 && 
b[18493] == 18493 && 
b[18494] == 18494 && 
b[18495] == 18495 && 
b[18496] == 18496 && 
b[18497] == 18497 && 
b[18498] == 18498 && 
b[18499] == 18499 && 
b[18500] == 18500 && 
b[18501] == 18501 && 
b[18502] == 18502 && 
b[18503] == 18503 && 
b[18504] == 18504 && 
b[18505] == 18505 && 
b[18506] == 18506 && 
b[18507] == 18507 && 
b[18508] == 18508 && 
b[18509] == 18509 && 
b[18510] == 18510 && 
b[18511] == 18511 && 
b[18512] == 18512 && 
b[18513] == 18513 && 
b[18514] == 18514 && 
b[18515] == 18515 && 
b[18516] == 18516 && 
b[18517] == 18517 && 
b[18518] == 18518 && 
b[18519] == 18519 && 
b[18520] == 18520 && 
b[18521] == 18521 && 
b[18522] == 18522 && 
b[18523] == 18523 && 
b[18524] == 18524 && 
b[18525] == 18525 && 
b[18526] == 18526 && 
b[18527] == 18527 && 
b[18528] == 18528 && 
b[18529] == 18529 && 
b[18530] == 18530 && 
b[18531] == 18531 && 
b[18532] == 18532 && 
b[18533] == 18533 && 
b[18534] == 18534 && 
b[18535] == 18535 && 
b[18536] == 18536 && 
b[18537] == 18537 && 
b[18538] == 18538 && 
b[18539] == 18539 && 
b[18540] == 18540 && 
b[18541] == 18541 && 
b[18542] == 18542 && 
b[18543] == 18543 && 
b[18544] == 18544 && 
b[18545] == 18545 && 
b[18546] == 18546 && 
b[18547] == 18547 && 
b[18548] == 18548 && 
b[18549] == 18549 && 
b[18550] == 18550 && 
b[18551] == 18551 && 
b[18552] == 18552 && 
b[18553] == 18553 && 
b[18554] == 18554 && 
b[18555] == 18555 && 
b[18556] == 18556 && 
b[18557] == 18557 && 
b[18558] == 18558 && 
b[18559] == 18559 && 
b[18560] == 18560 && 
b[18561] == 18561 && 
b[18562] == 18562 && 
b[18563] == 18563 && 
b[18564] == 18564 && 
b[18565] == 18565 && 
b[18566] == 18566 && 
b[18567] == 18567 && 
b[18568] == 18568 && 
b[18569] == 18569 && 
b[18570] == 18570 && 
b[18571] == 18571 && 
b[18572] == 18572 && 
b[18573] == 18573 && 
b[18574] == 18574 && 
b[18575] == 18575 && 
b[18576] == 18576 && 
b[18577] == 18577 && 
b[18578] == 18578 && 
b[18579] == 18579 && 
b[18580] == 18580 && 
b[18581] == 18581 && 
b[18582] == 18582 && 
b[18583] == 18583 && 
b[18584] == 18584 && 
b[18585] == 18585 && 
b[18586] == 18586 && 
b[18587] == 18587 && 
b[18588] == 18588 && 
b[18589] == 18589 && 
b[18590] == 18590 && 
b[18591] == 18591 && 
b[18592] == 18592 && 
b[18593] == 18593 && 
b[18594] == 18594 && 
b[18595] == 18595 && 
b[18596] == 18596 && 
b[18597] == 18597 && 
b[18598] == 18598 && 
b[18599] == 18599 && 
b[18600] == 18600 && 
b[18601] == 18601 && 
b[18602] == 18602 && 
b[18603] == 18603 && 
b[18604] == 18604 && 
b[18605] == 18605 && 
b[18606] == 18606 && 
b[18607] == 18607 && 
b[18608] == 18608 && 
b[18609] == 18609 && 
b[18610] == 18610 && 
b[18611] == 18611 && 
b[18612] == 18612 && 
b[18613] == 18613 && 
b[18614] == 18614 && 
b[18615] == 18615 && 
b[18616] == 18616 && 
b[18617] == 18617 && 
b[18618] == 18618 && 
b[18619] == 18619 && 
b[18620] == 18620 && 
b[18621] == 18621 && 
b[18622] == 18622 && 
b[18623] == 18623 && 
b[18624] == 18624 && 
b[18625] == 18625 && 
b[18626] == 18626 && 
b[18627] == 18627 && 
b[18628] == 18628 && 
b[18629] == 18629 && 
b[18630] == 18630 && 
b[18631] == 18631 && 
b[18632] == 18632 && 
b[18633] == 18633 && 
b[18634] == 18634 && 
b[18635] == 18635 && 
b[18636] == 18636 && 
b[18637] == 18637 && 
b[18638] == 18638 && 
b[18639] == 18639 && 
b[18640] == 18640 && 
b[18641] == 18641 && 
b[18642] == 18642 && 
b[18643] == 18643 && 
b[18644] == 18644 && 
b[18645] == 18645 && 
b[18646] == 18646 && 
b[18647] == 18647 && 
b[18648] == 18648 && 
b[18649] == 18649 && 
b[18650] == 18650 && 
b[18651] == 18651 && 
b[18652] == 18652 && 
b[18653] == 18653 && 
b[18654] == 18654 && 
b[18655] == 18655 && 
b[18656] == 18656 && 
b[18657] == 18657 && 
b[18658] == 18658 && 
b[18659] == 18659 && 
b[18660] == 18660 && 
b[18661] == 18661 && 
b[18662] == 18662 && 
b[18663] == 18663 && 
b[18664] == 18664 && 
b[18665] == 18665 && 
b[18666] == 18666 && 
b[18667] == 18667 && 
b[18668] == 18668 && 
b[18669] == 18669 && 
b[18670] == 18670 && 
b[18671] == 18671 && 
b[18672] == 18672 && 
b[18673] == 18673 && 
b[18674] == 18674 && 
b[18675] == 18675 && 
b[18676] == 18676 && 
b[18677] == 18677 && 
b[18678] == 18678 && 
b[18679] == 18679 && 
b[18680] == 18680 && 
b[18681] == 18681 && 
b[18682] == 18682 && 
b[18683] == 18683 && 
b[18684] == 18684 && 
b[18685] == 18685 && 
b[18686] == 18686 && 
b[18687] == 18687 && 
b[18688] == 18688 && 
b[18689] == 18689 && 
b[18690] == 18690 && 
b[18691] == 18691 && 
b[18692] == 18692 && 
b[18693] == 18693 && 
b[18694] == 18694 && 
b[18695] == 18695 && 
b[18696] == 18696 && 
b[18697] == 18697 && 
b[18698] == 18698 && 
b[18699] == 18699 && 
b[18700] == 18700 && 
b[18701] == 18701 && 
b[18702] == 18702 && 
b[18703] == 18703 && 
b[18704] == 18704 && 
b[18705] == 18705 && 
b[18706] == 18706 && 
b[18707] == 18707 && 
b[18708] == 18708 && 
b[18709] == 18709 && 
b[18710] == 18710 && 
b[18711] == 18711 && 
b[18712] == 18712 && 
b[18713] == 18713 && 
b[18714] == 18714 && 
b[18715] == 18715 && 
b[18716] == 18716 && 
b[18717] == 18717 && 
b[18718] == 18718 && 
b[18719] == 18719 && 
b[18720] == 18720 && 
b[18721] == 18721 && 
b[18722] == 18722 && 
b[18723] == 18723 && 
b[18724] == 18724 && 
b[18725] == 18725 && 
b[18726] == 18726 && 
b[18727] == 18727 && 
b[18728] == 18728 && 
b[18729] == 18729 && 
b[18730] == 18730 && 
b[18731] == 18731 && 
b[18732] == 18732 && 
b[18733] == 18733 && 
b[18734] == 18734 && 
b[18735] == 18735 && 
b[18736] == 18736 && 
b[18737] == 18737 && 
b[18738] == 18738 && 
b[18739] == 18739 && 
b[18740] == 18740 && 
b[18741] == 18741 && 
b[18742] == 18742 && 
b[18743] == 18743 && 
b[18744] == 18744 && 
b[18745] == 18745 && 
b[18746] == 18746 && 
b[18747] == 18747 && 
b[18748] == 18748 && 
b[18749] == 18749 && 
b[18750] == 18750 && 
b[18751] == 18751 && 
b[18752] == 18752 && 
b[18753] == 18753 && 
b[18754] == 18754 && 
b[18755] == 18755 && 
b[18756] == 18756 && 
b[18757] == 18757 && 
b[18758] == 18758 && 
b[18759] == 18759 && 
b[18760] == 18760 && 
b[18761] == 18761 && 
b[18762] == 18762 && 
b[18763] == 18763 && 
b[18764] == 18764 && 
b[18765] == 18765 && 
b[18766] == 18766 && 
b[18767] == 18767 && 
b[18768] == 18768 && 
b[18769] == 18769 && 
b[18770] == 18770 && 
b[18771] == 18771 && 
b[18772] == 18772 && 
b[18773] == 18773 && 
b[18774] == 18774 && 
b[18775] == 18775 && 
b[18776] == 18776 && 
b[18777] == 18777 && 
b[18778] == 18778 && 
b[18779] == 18779 && 
b[18780] == 18780 && 
b[18781] == 18781 && 
b[18782] == 18782 && 
b[18783] == 18783 && 
b[18784] == 18784 && 
b[18785] == 18785 && 
b[18786] == 18786 && 
b[18787] == 18787 && 
b[18788] == 18788 && 
b[18789] == 18789 && 
b[18790] == 18790 && 
b[18791] == 18791 && 
b[18792] == 18792 && 
b[18793] == 18793 && 
b[18794] == 18794 && 
b[18795] == 18795 && 
b[18796] == 18796 && 
b[18797] == 18797 && 
b[18798] == 18798 && 
b[18799] == 18799 && 
b[18800] == 18800 && 
b[18801] == 18801 && 
b[18802] == 18802 && 
b[18803] == 18803 && 
b[18804] == 18804 && 
b[18805] == 18805 && 
b[18806] == 18806 && 
b[18807] == 18807 && 
b[18808] == 18808 && 
b[18809] == 18809 && 
b[18810] == 18810 && 
b[18811] == 18811 && 
b[18812] == 18812 && 
b[18813] == 18813 && 
b[18814] == 18814 && 
b[18815] == 18815 && 
b[18816] == 18816 && 
b[18817] == 18817 && 
b[18818] == 18818 && 
b[18819] == 18819 && 
b[18820] == 18820 && 
b[18821] == 18821 && 
b[18822] == 18822 && 
b[18823] == 18823 && 
b[18824] == 18824 && 
b[18825] == 18825 && 
b[18826] == 18826 && 
b[18827] == 18827 && 
b[18828] == 18828 && 
b[18829] == 18829 && 
b[18830] == 18830 && 
b[18831] == 18831 && 
b[18832] == 18832 && 
b[18833] == 18833 && 
b[18834] == 18834 && 
b[18835] == 18835 && 
b[18836] == 18836 && 
b[18837] == 18837 && 
b[18838] == 18838 && 
b[18839] == 18839 && 
b[18840] == 18840 && 
b[18841] == 18841 && 
b[18842] == 18842 && 
b[18843] == 18843 && 
b[18844] == 18844 && 
b[18845] == 18845 && 
b[18846] == 18846 && 
b[18847] == 18847 && 
b[18848] == 18848 && 
b[18849] == 18849 && 
b[18850] == 18850 && 
b[18851] == 18851 && 
b[18852] == 18852 && 
b[18853] == 18853 && 
b[18854] == 18854 && 
b[18855] == 18855 && 
b[18856] == 18856 && 
b[18857] == 18857 && 
b[18858] == 18858 && 
b[18859] == 18859 && 
b[18860] == 18860 && 
b[18861] == 18861 && 
b[18862] == 18862 && 
b[18863] == 18863 && 
b[18864] == 18864 && 
b[18865] == 18865 && 
b[18866] == 18866 && 
b[18867] == 18867 && 
b[18868] == 18868 && 
b[18869] == 18869 && 
b[18870] == 18870 && 
b[18871] == 18871 && 
b[18872] == 18872 && 
b[18873] == 18873 && 
b[18874] == 18874 && 
b[18875] == 18875 && 
b[18876] == 18876 && 
b[18877] == 18877 && 
b[18878] == 18878 && 
b[18879] == 18879 && 
b[18880] == 18880 && 
b[18881] == 18881 && 
b[18882] == 18882 && 
b[18883] == 18883 && 
b[18884] == 18884 && 
b[18885] == 18885 && 
b[18886] == 18886 && 
b[18887] == 18887 && 
b[18888] == 18888 && 
b[18889] == 18889 && 
b[18890] == 18890 && 
b[18891] == 18891 && 
b[18892] == 18892 && 
b[18893] == 18893 && 
b[18894] == 18894 && 
b[18895] == 18895 && 
b[18896] == 18896 && 
b[18897] == 18897 && 
b[18898] == 18898 && 
b[18899] == 18899 && 
b[18900] == 18900 && 
b[18901] == 18901 && 
b[18902] == 18902 && 
b[18903] == 18903 && 
b[18904] == 18904 && 
b[18905] == 18905 && 
b[18906] == 18906 && 
b[18907] == 18907 && 
b[18908] == 18908 && 
b[18909] == 18909 && 
b[18910] == 18910 && 
b[18911] == 18911 && 
b[18912] == 18912 && 
b[18913] == 18913 && 
b[18914] == 18914 && 
b[18915] == 18915 && 
b[18916] == 18916 && 
b[18917] == 18917 && 
b[18918] == 18918 && 
b[18919] == 18919 && 
b[18920] == 18920 && 
b[18921] == 18921 && 
b[18922] == 18922 && 
b[18923] == 18923 && 
b[18924] == 18924 && 
b[18925] == 18925 && 
b[18926] == 18926 && 
b[18927] == 18927 && 
b[18928] == 18928 && 
b[18929] == 18929 && 
b[18930] == 18930 && 
b[18931] == 18931 && 
b[18932] == 18932 && 
b[18933] == 18933 && 
b[18934] == 18934 && 
b[18935] == 18935 && 
b[18936] == 18936 && 
b[18937] == 18937 && 
b[18938] == 18938 && 
b[18939] == 18939 && 
b[18940] == 18940 && 
b[18941] == 18941 && 
b[18942] == 18942 && 
b[18943] == 18943 && 
b[18944] == 18944 && 
b[18945] == 18945 && 
b[18946] == 18946 && 
b[18947] == 18947 && 
b[18948] == 18948 && 
b[18949] == 18949 && 
b[18950] == 18950 && 
b[18951] == 18951 && 
b[18952] == 18952 && 
b[18953] == 18953 && 
b[18954] == 18954 && 
b[18955] == 18955 && 
b[18956] == 18956 && 
b[18957] == 18957 && 
b[18958] == 18958 && 
b[18959] == 18959 && 
b[18960] == 18960 && 
b[18961] == 18961 && 
b[18962] == 18962 && 
b[18963] == 18963 && 
b[18964] == 18964 && 
b[18965] == 18965 && 
b[18966] == 18966 && 
b[18967] == 18967 && 
b[18968] == 18968 && 
b[18969] == 18969 && 
b[18970] == 18970 && 
b[18971] == 18971 && 
b[18972] == 18972 && 
b[18973] == 18973 && 
b[18974] == 18974 && 
b[18975] == 18975 && 
b[18976] == 18976 && 
b[18977] == 18977 && 
b[18978] == 18978 && 
b[18979] == 18979 && 
b[18980] == 18980 && 
b[18981] == 18981 && 
b[18982] == 18982 && 
b[18983] == 18983 && 
b[18984] == 18984 && 
b[18985] == 18985 && 
b[18986] == 18986 && 
b[18987] == 18987 && 
b[18988] == 18988 && 
b[18989] == 18989 && 
b[18990] == 18990 && 
b[18991] == 18991 && 
b[18992] == 18992 && 
b[18993] == 18993 && 
b[18994] == 18994 && 
b[18995] == 18995 && 
b[18996] == 18996 && 
b[18997] == 18997 && 
b[18998] == 18998 && 
b[18999] == 18999 && 
b[19000] == 19000 && 
b[19001] == 19001 && 
b[19002] == 19002 && 
b[19003] == 19003 && 
b[19004] == 19004 && 
b[19005] == 19005 && 
b[19006] == 19006 && 
b[19007] == 19007 && 
b[19008] == 19008 && 
b[19009] == 19009 && 
b[19010] == 19010 && 
b[19011] == 19011 && 
b[19012] == 19012 && 
b[19013] == 19013 && 
b[19014] == 19014 && 
b[19015] == 19015 && 
b[19016] == 19016 && 
b[19017] == 19017 && 
b[19018] == 19018 && 
b[19019] == 19019 && 
b[19020] == 19020 && 
b[19021] == 19021 && 
b[19022] == 19022 && 
b[19023] == 19023 && 
b[19024] == 19024 && 
b[19025] == 19025 && 
b[19026] == 19026 && 
b[19027] == 19027 && 
b[19028] == 19028 && 
b[19029] == 19029 && 
b[19030] == 19030 && 
b[19031] == 19031 && 
b[19032] == 19032 && 
b[19033] == 19033 && 
b[19034] == 19034 && 
b[19035] == 19035 && 
b[19036] == 19036 && 
b[19037] == 19037 && 
b[19038] == 19038 && 
b[19039] == 19039 && 
b[19040] == 19040 && 
b[19041] == 19041 && 
b[19042] == 19042 && 
b[19043] == 19043 && 
b[19044] == 19044 && 
b[19045] == 19045 && 
b[19046] == 19046 && 
b[19047] == 19047 && 
b[19048] == 19048 && 
b[19049] == 19049 && 
b[19050] == 19050 && 
b[19051] == 19051 && 
b[19052] == 19052 && 
b[19053] == 19053 && 
b[19054] == 19054 && 
b[19055] == 19055 && 
b[19056] == 19056 && 
b[19057] == 19057 && 
b[19058] == 19058 && 
b[19059] == 19059 && 
b[19060] == 19060 && 
b[19061] == 19061 && 
b[19062] == 19062 && 
b[19063] == 19063 && 
b[19064] == 19064 && 
b[19065] == 19065 && 
b[19066] == 19066 && 
b[19067] == 19067 && 
b[19068] == 19068 && 
b[19069] == 19069 && 
b[19070] == 19070 && 
b[19071] == 19071 && 
b[19072] == 19072 && 
b[19073] == 19073 && 
b[19074] == 19074 && 
b[19075] == 19075 && 
b[19076] == 19076 && 
b[19077] == 19077 && 
b[19078] == 19078 && 
b[19079] == 19079 && 
b[19080] == 19080 && 
b[19081] == 19081 && 
b[19082] == 19082 && 
b[19083] == 19083 && 
b[19084] == 19084 && 
b[19085] == 19085 && 
b[19086] == 19086 && 
b[19087] == 19087 && 
b[19088] == 19088 && 
b[19089] == 19089 && 
b[19090] == 19090 && 
b[19091] == 19091 && 
b[19092] == 19092 && 
b[19093] == 19093 && 
b[19094] == 19094 && 
b[19095] == 19095 && 
b[19096] == 19096 && 
b[19097] == 19097 && 
b[19098] == 19098 && 
b[19099] == 19099 && 
b[19100] == 19100 && 
b[19101] == 19101 && 
b[19102] == 19102 && 
b[19103] == 19103 && 
b[19104] == 19104 && 
b[19105] == 19105 && 
b[19106] == 19106 && 
b[19107] == 19107 && 
b[19108] == 19108 && 
b[19109] == 19109 && 
b[19110] == 19110 && 
b[19111] == 19111 && 
b[19112] == 19112 && 
b[19113] == 19113 && 
b[19114] == 19114 && 
b[19115] == 19115 && 
b[19116] == 19116 && 
b[19117] == 19117 && 
b[19118] == 19118 && 
b[19119] == 19119 && 
b[19120] == 19120 && 
b[19121] == 19121 && 
b[19122] == 19122 && 
b[19123] == 19123 && 
b[19124] == 19124 && 
b[19125] == 19125 && 
b[19126] == 19126 && 
b[19127] == 19127 && 
b[19128] == 19128 && 
b[19129] == 19129 && 
b[19130] == 19130 && 
b[19131] == 19131 && 
b[19132] == 19132 && 
b[19133] == 19133 && 
b[19134] == 19134 && 
b[19135] == 19135 && 
b[19136] == 19136 && 
b[19137] == 19137 && 
b[19138] == 19138 && 
b[19139] == 19139 && 
b[19140] == 19140 && 
b[19141] == 19141 && 
b[19142] == 19142 && 
b[19143] == 19143 && 
b[19144] == 19144 && 
b[19145] == 19145 && 
b[19146] == 19146 && 
b[19147] == 19147 && 
b[19148] == 19148 && 
b[19149] == 19149 && 
b[19150] == 19150 && 
b[19151] == 19151 && 
b[19152] == 19152 && 
b[19153] == 19153 && 
b[19154] == 19154 && 
b[19155] == 19155 && 
b[19156] == 19156 && 
b[19157] == 19157 && 
b[19158] == 19158 && 
b[19159] == 19159 && 
b[19160] == 19160 && 
b[19161] == 19161 && 
b[19162] == 19162 && 
b[19163] == 19163 && 
b[19164] == 19164 && 
b[19165] == 19165 && 
b[19166] == 19166 && 
b[19167] == 19167 && 
b[19168] == 19168 && 
b[19169] == 19169 && 
b[19170] == 19170 && 
b[19171] == 19171 && 
b[19172] == 19172 && 
b[19173] == 19173 && 
b[19174] == 19174 && 
b[19175] == 19175 && 
b[19176] == 19176 && 
b[19177] == 19177 && 
b[19178] == 19178 && 
b[19179] == 19179 && 
b[19180] == 19180 && 
b[19181] == 19181 && 
b[19182] == 19182 && 
b[19183] == 19183 && 
b[19184] == 19184 && 
b[19185] == 19185 && 
b[19186] == 19186 && 
b[19187] == 19187 && 
b[19188] == 19188 && 
b[19189] == 19189 && 
b[19190] == 19190 && 
b[19191] == 19191 && 
b[19192] == 19192 && 
b[19193] == 19193 && 
b[19194] == 19194 && 
b[19195] == 19195 && 
b[19196] == 19196 && 
b[19197] == 19197 && 
b[19198] == 19198 && 
b[19199] == 19199 && 
b[19200] == 19200 && 
b[19201] == 19201 && 
b[19202] == 19202 && 
b[19203] == 19203 && 
b[19204] == 19204 && 
b[19205] == 19205 && 
b[19206] == 19206 && 
b[19207] == 19207 && 
b[19208] == 19208 && 
b[19209] == 19209 && 
b[19210] == 19210 && 
b[19211] == 19211 && 
b[19212] == 19212 && 
b[19213] == 19213 && 
b[19214] == 19214 && 
b[19215] == 19215 && 
b[19216] == 19216 && 
b[19217] == 19217 && 
b[19218] == 19218 && 
b[19219] == 19219 && 
b[19220] == 19220 && 
b[19221] == 19221 && 
b[19222] == 19222 && 
b[19223] == 19223 && 
b[19224] == 19224 && 
b[19225] == 19225 && 
b[19226] == 19226 && 
b[19227] == 19227 && 
b[19228] == 19228 && 
b[19229] == 19229 && 
b[19230] == 19230 && 
b[19231] == 19231 && 
b[19232] == 19232 && 
b[19233] == 19233 && 
b[19234] == 19234 && 
b[19235] == 19235 && 
b[19236] == 19236 && 
b[19237] == 19237 && 
b[19238] == 19238 && 
b[19239] == 19239 && 
b[19240] == 19240 && 
b[19241] == 19241 && 
b[19242] == 19242 && 
b[19243] == 19243 && 
b[19244] == 19244 && 
b[19245] == 19245 && 
b[19246] == 19246 && 
b[19247] == 19247 && 
b[19248] == 19248 && 
b[19249] == 19249 && 
b[19250] == 19250 && 
b[19251] == 19251 && 
b[19252] == 19252 && 
b[19253] == 19253 && 
b[19254] == 19254 && 
b[19255] == 19255 && 
b[19256] == 19256 && 
b[19257] == 19257 && 
b[19258] == 19258 && 
b[19259] == 19259 && 
b[19260] == 19260 && 
b[19261] == 19261 && 
b[19262] == 19262 && 
b[19263] == 19263 && 
b[19264] == 19264 && 
b[19265] == 19265 && 
b[19266] == 19266 && 
b[19267] == 19267 && 
b[19268] == 19268 && 
b[19269] == 19269 && 
b[19270] == 19270 && 
b[19271] == 19271 && 
b[19272] == 19272 && 
b[19273] == 19273 && 
b[19274] == 19274 && 
b[19275] == 19275 && 
b[19276] == 19276 && 
b[19277] == 19277 && 
b[19278] == 19278 && 
b[19279] == 19279 && 
b[19280] == 19280 && 
b[19281] == 19281 && 
b[19282] == 19282 && 
b[19283] == 19283 && 
b[19284] == 19284 && 
b[19285] == 19285 && 
b[19286] == 19286 && 
b[19287] == 19287 && 
b[19288] == 19288 && 
b[19289] == 19289 && 
b[19290] == 19290 && 
b[19291] == 19291 && 
b[19292] == 19292 && 
b[19293] == 19293 && 
b[19294] == 19294 && 
b[19295] == 19295 && 
b[19296] == 19296 && 
b[19297] == 19297 && 
b[19298] == 19298 && 
b[19299] == 19299 && 
b[19300] == 19300 && 
b[19301] == 19301 && 
b[19302] == 19302 && 
b[19303] == 19303 && 
b[19304] == 19304 && 
b[19305] == 19305 && 
b[19306] == 19306 && 
b[19307] == 19307 && 
b[19308] == 19308 && 
b[19309] == 19309 && 
b[19310] == 19310 && 
b[19311] == 19311 && 
b[19312] == 19312 && 
b[19313] == 19313 && 
b[19314] == 19314 && 
b[19315] == 19315 && 
b[19316] == 19316 && 
b[19317] == 19317 && 
b[19318] == 19318 && 
b[19319] == 19319 && 
b[19320] == 19320 && 
b[19321] == 19321 && 
b[19322] == 19322 && 
b[19323] == 19323 && 
b[19324] == 19324 && 
b[19325] == 19325 && 
b[19326] == 19326 && 
b[19327] == 19327 && 
b[19328] == 19328 && 
b[19329] == 19329 && 
b[19330] == 19330 && 
b[19331] == 19331 && 
b[19332] == 19332 && 
b[19333] == 19333 && 
b[19334] == 19334 && 
b[19335] == 19335 && 
b[19336] == 19336 && 
b[19337] == 19337 && 
b[19338] == 19338 && 
b[19339] == 19339 && 
b[19340] == 19340 && 
b[19341] == 19341 && 
b[19342] == 19342 && 
b[19343] == 19343 && 
b[19344] == 19344 && 
b[19345] == 19345 && 
b[19346] == 19346 && 
b[19347] == 19347 && 
b[19348] == 19348 && 
b[19349] == 19349 && 
b[19350] == 19350 && 
b[19351] == 19351 && 
b[19352] == 19352 && 
b[19353] == 19353 && 
b[19354] == 19354 && 
b[19355] == 19355 && 
b[19356] == 19356 && 
b[19357] == 19357 && 
b[19358] == 19358 && 
b[19359] == 19359 && 
b[19360] == 19360 && 
b[19361] == 19361 && 
b[19362] == 19362 && 
b[19363] == 19363 && 
b[19364] == 19364 && 
b[19365] == 19365 && 
b[19366] == 19366 && 
b[19367] == 19367 && 
b[19368] == 19368 && 
b[19369] == 19369 && 
b[19370] == 19370 && 
b[19371] == 19371 && 
b[19372] == 19372 && 
b[19373] == 19373 && 
b[19374] == 19374 && 
b[19375] == 19375 && 
b[19376] == 19376 && 
b[19377] == 19377 && 
b[19378] == 19378 && 
b[19379] == 19379 && 
b[19380] == 19380 && 
b[19381] == 19381 && 
b[19382] == 19382 && 
b[19383] == 19383 && 
b[19384] == 19384 && 
b[19385] == 19385 && 
b[19386] == 19386 && 
b[19387] == 19387 && 
b[19388] == 19388 && 
b[19389] == 19389 && 
b[19390] == 19390 && 
b[19391] == 19391 && 
b[19392] == 19392 && 
b[19393] == 19393 && 
b[19394] == 19394 && 
b[19395] == 19395 && 
b[19396] == 19396 && 
b[19397] == 19397 && 
b[19398] == 19398 && 
b[19399] == 19399 && 
b[19400] == 19400 && 
b[19401] == 19401 && 
b[19402] == 19402 && 
b[19403] == 19403 && 
b[19404] == 19404 && 
b[19405] == 19405 && 
b[19406] == 19406 && 
b[19407] == 19407 && 
b[19408] == 19408 && 
b[19409] == 19409 && 
b[19410] == 19410 && 
b[19411] == 19411 && 
b[19412] == 19412 && 
b[19413] == 19413 && 
b[19414] == 19414 && 
b[19415] == 19415 && 
b[19416] == 19416 && 
b[19417] == 19417 && 
b[19418] == 19418 && 
b[19419] == 19419 && 
b[19420] == 19420 && 
b[19421] == 19421 && 
b[19422] == 19422 && 
b[19423] == 19423 && 
b[19424] == 19424 && 
b[19425] == 19425 && 
b[19426] == 19426 && 
b[19427] == 19427 && 
b[19428] == 19428 && 
b[19429] == 19429 && 
b[19430] == 19430 && 
b[19431] == 19431 && 
b[19432] == 19432 && 
b[19433] == 19433 && 
b[19434] == 19434 && 
b[19435] == 19435 && 
b[19436] == 19436 && 
b[19437] == 19437 && 
b[19438] == 19438 && 
b[19439] == 19439 && 
b[19440] == 19440 && 
b[19441] == 19441 && 
b[19442] == 19442 && 
b[19443] == 19443 && 
b[19444] == 19444 && 
b[19445] == 19445 && 
b[19446] == 19446 && 
b[19447] == 19447 && 
b[19448] == 19448 && 
b[19449] == 19449 && 
b[19450] == 19450 && 
b[19451] == 19451 && 
b[19452] == 19452 && 
b[19453] == 19453 && 
b[19454] == 19454 && 
b[19455] == 19455 && 
b[19456] == 19456 && 
b[19457] == 19457 && 
b[19458] == 19458 && 
b[19459] == 19459 && 
b[19460] == 19460 && 
b[19461] == 19461 && 
b[19462] == 19462 && 
b[19463] == 19463 && 
b[19464] == 19464 && 
b[19465] == 19465 && 
b[19466] == 19466 && 
b[19467] == 19467 && 
b[19468] == 19468 && 
b[19469] == 19469 && 
b[19470] == 19470 && 
b[19471] == 19471 && 
b[19472] == 19472 && 
b[19473] == 19473 && 
b[19474] == 19474 && 
b[19475] == 19475 && 
b[19476] == 19476 && 
b[19477] == 19477 && 
b[19478] == 19478 && 
b[19479] == 19479 && 
b[19480] == 19480 && 
b[19481] == 19481 && 
b[19482] == 19482 && 
b[19483] == 19483 && 
b[19484] == 19484 && 
b[19485] == 19485 && 
b[19486] == 19486 && 
b[19487] == 19487 && 
b[19488] == 19488 && 
b[19489] == 19489 && 
b[19490] == 19490 && 
b[19491] == 19491 && 
b[19492] == 19492 && 
b[19493] == 19493 && 
b[19494] == 19494 && 
b[19495] == 19495 && 
b[19496] == 19496 && 
b[19497] == 19497 && 
b[19498] == 19498 && 
b[19499] == 19499 && 
b[19500] == 19500 && 
b[19501] == 19501 && 
b[19502] == 19502 && 
b[19503] == 19503 && 
b[19504] == 19504 && 
b[19505] == 19505 && 
b[19506] == 19506 && 
b[19507] == 19507 && 
b[19508] == 19508 && 
b[19509] == 19509 && 
b[19510] == 19510 && 
b[19511] == 19511 && 
b[19512] == 19512 && 
b[19513] == 19513 && 
b[19514] == 19514 && 
b[19515] == 19515 && 
b[19516] == 19516 && 
b[19517] == 19517 && 
b[19518] == 19518 && 
b[19519] == 19519 && 
b[19520] == 19520 && 
b[19521] == 19521 && 
b[19522] == 19522 && 
b[19523] == 19523 && 
b[19524] == 19524 && 
b[19525] == 19525 && 
b[19526] == 19526 && 
b[19527] == 19527 && 
b[19528] == 19528 && 
b[19529] == 19529 && 
b[19530] == 19530 && 
b[19531] == 19531 && 
b[19532] == 19532 && 
b[19533] == 19533 && 
b[19534] == 19534 && 
b[19535] == 19535 && 
b[19536] == 19536 && 
b[19537] == 19537 && 
b[19538] == 19538 && 
b[19539] == 19539 && 
b[19540] == 19540 && 
b[19541] == 19541 && 
b[19542] == 19542 && 
b[19543] == 19543 && 
b[19544] == 19544 && 
b[19545] == 19545 && 
b[19546] == 19546 && 
b[19547] == 19547 && 
b[19548] == 19548 && 
b[19549] == 19549 && 
b[19550] == 19550 && 
b[19551] == 19551 && 
b[19552] == 19552 && 
b[19553] == 19553 && 
b[19554] == 19554 && 
b[19555] == 19555 && 
b[19556] == 19556 && 
b[19557] == 19557 && 
b[19558] == 19558 && 
b[19559] == 19559 && 
b[19560] == 19560 && 
b[19561] == 19561 && 
b[19562] == 19562 && 
b[19563] == 19563 && 
b[19564] == 19564 && 
b[19565] == 19565 && 
b[19566] == 19566 && 
b[19567] == 19567 && 
b[19568] == 19568 && 
b[19569] == 19569 && 
b[19570] == 19570 && 
b[19571] == 19571 && 
b[19572] == 19572 && 
b[19573] == 19573 && 
b[19574] == 19574 && 
b[19575] == 19575 && 
b[19576] == 19576 && 
b[19577] == 19577 && 
b[19578] == 19578 && 
b[19579] == 19579 && 
b[19580] == 19580 && 
b[19581] == 19581 && 
b[19582] == 19582 && 
b[19583] == 19583 && 
b[19584] == 19584 && 
b[19585] == 19585 && 
b[19586] == 19586 && 
b[19587] == 19587 && 
b[19588] == 19588 && 
b[19589] == 19589 && 
b[19590] == 19590 && 
b[19591] == 19591 && 
b[19592] == 19592 && 
b[19593] == 19593 && 
b[19594] == 19594 && 
b[19595] == 19595 && 
b[19596] == 19596 && 
b[19597] == 19597 && 
b[19598] == 19598 && 
b[19599] == 19599 && 
b[19600] == 19600 && 
b[19601] == 19601 && 
b[19602] == 19602 && 
b[19603] == 19603 && 
b[19604] == 19604 && 
b[19605] == 19605 && 
b[19606] == 19606 && 
b[19607] == 19607 && 
b[19608] == 19608 && 
b[19609] == 19609 && 
b[19610] == 19610 && 
b[19611] == 19611 && 
b[19612] == 19612 && 
b[19613] == 19613 && 
b[19614] == 19614 && 
b[19615] == 19615 && 
b[19616] == 19616 && 
b[19617] == 19617 && 
b[19618] == 19618 && 
b[19619] == 19619 && 
b[19620] == 19620 && 
b[19621] == 19621 && 
b[19622] == 19622 && 
b[19623] == 19623 && 
b[19624] == 19624 && 
b[19625] == 19625 && 
b[19626] == 19626 && 
b[19627] == 19627 && 
b[19628] == 19628 && 
b[19629] == 19629 && 
b[19630] == 19630 && 
b[19631] == 19631 && 
b[19632] == 19632 && 
b[19633] == 19633 && 
b[19634] == 19634 && 
b[19635] == 19635 && 
b[19636] == 19636 && 
b[19637] == 19637 && 
b[19638] == 19638 && 
b[19639] == 19639 && 
b[19640] == 19640 && 
b[19641] == 19641 && 
b[19642] == 19642 && 
b[19643] == 19643 && 
b[19644] == 19644 && 
b[19645] == 19645 && 
b[19646] == 19646 && 
b[19647] == 19647 && 
b[19648] == 19648 && 
b[19649] == 19649 && 
b[19650] == 19650 && 
b[19651] == 19651 && 
b[19652] == 19652 && 
b[19653] == 19653 && 
b[19654] == 19654 && 
b[19655] == 19655 && 
b[19656] == 19656 && 
b[19657] == 19657 && 
b[19658] == 19658 && 
b[19659] == 19659 && 
b[19660] == 19660 && 
b[19661] == 19661 && 
b[19662] == 19662 && 
b[19663] == 19663 && 
b[19664] == 19664 && 
b[19665] == 19665 && 
b[19666] == 19666 && 
b[19667] == 19667 && 
b[19668] == 19668 && 
b[19669] == 19669 && 
b[19670] == 19670 && 
b[19671] == 19671 && 
b[19672] == 19672 && 
b[19673] == 19673 && 
b[19674] == 19674 && 
b[19675] == 19675 && 
b[19676] == 19676 && 
b[19677] == 19677 && 
b[19678] == 19678 && 
b[19679] == 19679 && 
b[19680] == 19680 && 
b[19681] == 19681 && 
b[19682] == 19682 && 
b[19683] == 19683 && 
b[19684] == 19684 && 
b[19685] == 19685 && 
b[19686] == 19686 && 
b[19687] == 19687 && 
b[19688] == 19688 && 
b[19689] == 19689 && 
b[19690] == 19690 && 
b[19691] == 19691 && 
b[19692] == 19692 && 
b[19693] == 19693 && 
b[19694] == 19694 && 
b[19695] == 19695 && 
b[19696] == 19696 && 
b[19697] == 19697 && 
b[19698] == 19698 && 
b[19699] == 19699 && 
b[19700] == 19700 && 
b[19701] == 19701 && 
b[19702] == 19702 && 
b[19703] == 19703 && 
b[19704] == 19704 && 
b[19705] == 19705 && 
b[19706] == 19706 && 
b[19707] == 19707 && 
b[19708] == 19708 && 
b[19709] == 19709 && 
b[19710] == 19710 && 
b[19711] == 19711 && 
b[19712] == 19712 && 
b[19713] == 19713 && 
b[19714] == 19714 && 
b[19715] == 19715 && 
b[19716] == 19716 && 
b[19717] == 19717 && 
b[19718] == 19718 && 
b[19719] == 19719 && 
b[19720] == 19720 && 
b[19721] == 19721 && 
b[19722] == 19722 && 
b[19723] == 19723 && 
b[19724] == 19724 && 
b[19725] == 19725 && 
b[19726] == 19726 && 
b[19727] == 19727 && 
b[19728] == 19728 && 
b[19729] == 19729 && 
b[19730] == 19730 && 
b[19731] == 19731 && 
b[19732] == 19732 && 
b[19733] == 19733 && 
b[19734] == 19734 && 
b[19735] == 19735 && 
b[19736] == 19736 && 
b[19737] == 19737 && 
b[19738] == 19738 && 
b[19739] == 19739 && 
b[19740] == 19740 && 
b[19741] == 19741 && 
b[19742] == 19742 && 
b[19743] == 19743 && 
b[19744] == 19744 && 
b[19745] == 19745 && 
b[19746] == 19746 && 
b[19747] == 19747 && 
b[19748] == 19748 && 
b[19749] == 19749 && 
b[19750] == 19750 && 
b[19751] == 19751 && 
b[19752] == 19752 && 
b[19753] == 19753 && 
b[19754] == 19754 && 
b[19755] == 19755 && 
b[19756] == 19756 && 
b[19757] == 19757 && 
b[19758] == 19758 && 
b[19759] == 19759 && 
b[19760] == 19760 && 
b[19761] == 19761 && 
b[19762] == 19762 && 
b[19763] == 19763 && 
b[19764] == 19764 && 
b[19765] == 19765 && 
b[19766] == 19766 && 
b[19767] == 19767 && 
b[19768] == 19768 && 
b[19769] == 19769 && 
b[19770] == 19770 && 
b[19771] == 19771 && 
b[19772] == 19772 && 
b[19773] == 19773 && 
b[19774] == 19774 && 
b[19775] == 19775 && 
b[19776] == 19776 && 
b[19777] == 19777 && 
b[19778] == 19778 && 
b[19779] == 19779 && 
b[19780] == 19780 && 
b[19781] == 19781 && 
b[19782] == 19782 && 
b[19783] == 19783 && 
b[19784] == 19784 && 
b[19785] == 19785 && 
b[19786] == 19786 && 
b[19787] == 19787 && 
b[19788] == 19788 && 
b[19789] == 19789 && 
b[19790] == 19790 && 
b[19791] == 19791 && 
b[19792] == 19792 && 
b[19793] == 19793 && 
b[19794] == 19794 && 
b[19795] == 19795 && 
b[19796] == 19796 && 
b[19797] == 19797 && 
b[19798] == 19798 && 
b[19799] == 19799 && 
b[19800] == 19800 && 
b[19801] == 19801 && 
b[19802] == 19802 && 
b[19803] == 19803 && 
b[19804] == 19804 && 
b[19805] == 19805 && 
b[19806] == 19806 && 
b[19807] == 19807 && 
b[19808] == 19808 && 
b[19809] == 19809 && 
b[19810] == 19810 && 
b[19811] == 19811 && 
b[19812] == 19812 && 
b[19813] == 19813 && 
b[19814] == 19814 && 
b[19815] == 19815 && 
b[19816] == 19816 && 
b[19817] == 19817 && 
b[19818] == 19818 && 
b[19819] == 19819 && 
b[19820] == 19820 && 
b[19821] == 19821 && 
b[19822] == 19822 && 
b[19823] == 19823 && 
b[19824] == 19824 && 
b[19825] == 19825 && 
b[19826] == 19826 && 
b[19827] == 19827 && 
b[19828] == 19828 && 
b[19829] == 19829 && 
b[19830] == 19830 && 
b[19831] == 19831 && 
b[19832] == 19832 && 
b[19833] == 19833 && 
b[19834] == 19834 && 
b[19835] == 19835 && 
b[19836] == 19836 && 
b[19837] == 19837 && 
b[19838] == 19838 && 
b[19839] == 19839 && 
b[19840] == 19840 && 
b[19841] == 19841 && 
b[19842] == 19842 && 
b[19843] == 19843 && 
b[19844] == 19844 && 
b[19845] == 19845 && 
b[19846] == 19846 && 
b[19847] == 19847 && 
b[19848] == 19848 && 
b[19849] == 19849 && 
b[19850] == 19850 && 
b[19851] == 19851 && 
b[19852] == 19852 && 
b[19853] == 19853 && 
b[19854] == 19854 && 
b[19855] == 19855 && 
b[19856] == 19856 && 
b[19857] == 19857 && 
b[19858] == 19858 && 
b[19859] == 19859 && 
b[19860] == 19860 && 
b[19861] == 19861 && 
b[19862] == 19862 && 
b[19863] == 19863 && 
b[19864] == 19864 && 
b[19865] == 19865 && 
b[19866] == 19866 && 
b[19867] == 19867 && 
b[19868] == 19868 && 
b[19869] == 19869 && 
b[19870] == 19870 && 
b[19871] == 19871 && 
b[19872] == 19872 && 
b[19873] == 19873 && 
b[19874] == 19874 && 
b[19875] == 19875 && 
b[19876] == 19876 && 
b[19877] == 19877 && 
b[19878] == 19878 && 
b[19879] == 19879 && 
b[19880] == 19880 && 
b[19881] == 19881 && 
b[19882] == 19882 && 
b[19883] == 19883 && 
b[19884] == 19884 && 
b[19885] == 19885 && 
b[19886] == 19886 && 
b[19887] == 19887 && 
b[19888] == 19888 && 
b[19889] == 19889 && 
b[19890] == 19890 && 
b[19891] == 19891 && 
b[19892] == 19892 && 
b[19893] == 19893 && 
b[19894] == 19894 && 
b[19895] == 19895 && 
b[19896] == 19896 && 
b[19897] == 19897 && 
b[19898] == 19898 && 
b[19899] == 19899 && 
b[19900] == 19900 && 
b[19901] == 19901 && 
b[19902] == 19902 && 
b[19903] == 19903 && 
b[19904] == 19904 && 
b[19905] == 19905 && 
b[19906] == 19906 && 
b[19907] == 19907 && 
b[19908] == 19908 && 
b[19909] == 19909 && 
b[19910] == 19910 && 
b[19911] == 19911 && 
b[19912] == 19912 && 
b[19913] == 19913 && 
b[19914] == 19914 && 
b[19915] == 19915 && 
b[19916] == 19916 && 
b[19917] == 19917 && 
b[19918] == 19918 && 
b[19919] == 19919 && 
b[19920] == 19920 && 
b[19921] == 19921 && 
b[19922] == 19922 && 
b[19923] == 19923 && 
b[19924] == 19924 && 
b[19925] == 19925 && 
b[19926] == 19926 && 
b[19927] == 19927 && 
b[19928] == 19928 && 
b[19929] == 19929 && 
b[19930] == 19930 && 
b[19931] == 19931 && 
b[19932] == 19932 && 
b[19933] == 19933 && 
b[19934] == 19934 && 
b[19935] == 19935 && 
b[19936] == 19936 && 
b[19937] == 19937 && 
b[19938] == 19938 && 
b[19939] == 19939 && 
b[19940] == 19940 && 
b[19941] == 19941 && 
b[19942] == 19942 && 
b[19943] == 19943 && 
b[19944] == 19944 && 
b[19945] == 19945 && 
b[19946] == 19946 && 
b[19947] == 19947 && 
b[19948] == 19948 && 
b[19949] == 19949 && 
b[19950] == 19950 && 
b[19951] == 19951 && 
b[19952] == 19952 && 
b[19953] == 19953 && 
b[19954] == 19954 && 
b[19955] == 19955 && 
b[19956] == 19956 && 
b[19957] == 19957 && 
b[19958] == 19958 && 
b[19959] == 19959 && 
b[19960] == 19960 && 
b[19961] == 19961 && 
b[19962] == 19962 && 
b[19963] == 19963 && 
b[19964] == 19964 && 
b[19965] == 19965 && 
b[19966] == 19966 && 
b[19967] == 19967 && 
b[19968] == 19968 && 
b[19969] == 19969 && 
b[19970] == 19970 && 
b[19971] == 19971 && 
b[19972] == 19972 && 
b[19973] == 19973 && 
b[19974] == 19974 && 
b[19975] == 19975 && 
b[19976] == 19976 && 
b[19977] == 19977 && 
b[19978] == 19978 && 
b[19979] == 19979 && 
b[19980] == 19980 && 
b[19981] == 19981 && 
b[19982] == 19982 && 
b[19983] == 19983 && 
b[19984] == 19984 && 
b[19985] == 19985 && 
b[19986] == 19986 && 
b[19987] == 19987 && 
b[19988] == 19988 && 
b[19989] == 19989 && 
b[19990] == 19990 && 
b[19991] == 19991 && 
b[19992] == 19992 && 
b[19993] == 19993 && 
b[19994] == 19994 && 
b[19995] == 19995 && 
b[19996] == 19996 && 
b[19997] == 19997 && 
b[19998] == 19998 && 
b[19999] == 19999 && 
b[20000] == 20000 && 
b[20001] == 20001 && 
b[20002] == 20002 && 
b[20003] == 20003 && 
b[20004] == 20004 && 
b[20005] == 20005 && 
b[20006] == 20006 && 
b[20007] == 20007 && 
b[20008] == 20008 && 
b[20009] == 20009 && 
b[20010] == 20010 && 
b[20011] == 20011 && 
b[20012] == 20012 && 
b[20013] == 20013 && 
b[20014] == 20014 && 
b[20015] == 20015 && 
b[20016] == 20016 && 
b[20017] == 20017 && 
b[20018] == 20018 && 
b[20019] == 20019 && 
b[20020] == 20020 && 
b[20021] == 20021 && 
b[20022] == 20022 && 
b[20023] == 20023 && 
b[20024] == 20024 && 
b[20025] == 20025 && 
b[20026] == 20026 && 
b[20027] == 20027 && 
b[20028] == 20028 && 
b[20029] == 20029 && 
b[20030] == 20030 && 
b[20031] == 20031 && 
b[20032] == 20032 && 
b[20033] == 20033 && 
b[20034] == 20034 && 
b[20035] == 20035 && 
b[20036] == 20036 && 
b[20037] == 20037 && 
b[20038] == 20038 && 
b[20039] == 20039 && 
b[20040] == 20040 && 
b[20041] == 20041 && 
b[20042] == 20042 && 
b[20043] == 20043 && 
b[20044] == 20044 && 
b[20045] == 20045 && 
b[20046] == 20046 && 
b[20047] == 20047 && 
b[20048] == 20048 && 
b[20049] == 20049 && 
b[20050] == 20050 && 
b[20051] == 20051 && 
b[20052] == 20052 && 
b[20053] == 20053 && 
b[20054] == 20054 && 
b[20055] == 20055 && 
b[20056] == 20056 && 
b[20057] == 20057 && 
b[20058] == 20058 && 
b[20059] == 20059 && 
b[20060] == 20060 && 
b[20061] == 20061 && 
b[20062] == 20062 && 
b[20063] == 20063 && 
b[20064] == 20064 && 
b[20065] == 20065 && 
b[20066] == 20066 && 
b[20067] == 20067 && 
b[20068] == 20068 && 
b[20069] == 20069 && 
b[20070] == 20070 && 
b[20071] == 20071 && 
b[20072] == 20072 && 
b[20073] == 20073 && 
b[20074] == 20074 && 
b[20075] == 20075 && 
b[20076] == 20076 && 
b[20077] == 20077 && 
b[20078] == 20078 && 
b[20079] == 20079 && 
b[20080] == 20080 && 
b[20081] == 20081 && 
b[20082] == 20082 && 
b[20083] == 20083 && 
b[20084] == 20084 && 
b[20085] == 20085 && 
b[20086] == 20086 && 
b[20087] == 20087 && 
b[20088] == 20088 && 
b[20089] == 20089 && 
b[20090] == 20090 && 
b[20091] == 20091 && 
b[20092] == 20092 && 
b[20093] == 20093 && 
b[20094] == 20094 && 
b[20095] == 20095 && 
b[20096] == 20096 && 
b[20097] == 20097 && 
b[20098] == 20098 && 
b[20099] == 20099 && 
b[20100] == 20100 && 
b[20101] == 20101 && 
b[20102] == 20102 && 
b[20103] == 20103 && 
b[20104] == 20104 && 
b[20105] == 20105 && 
b[20106] == 20106 && 
b[20107] == 20107 && 
b[20108] == 20108 && 
b[20109] == 20109 && 
b[20110] == 20110 && 
b[20111] == 20111 && 
b[20112] == 20112 && 
b[20113] == 20113 && 
b[20114] == 20114 && 
b[20115] == 20115 && 
b[20116] == 20116 && 
b[20117] == 20117 && 
b[20118] == 20118 && 
b[20119] == 20119 && 
b[20120] == 20120 && 
b[20121] == 20121 && 
b[20122] == 20122 && 
b[20123] == 20123 && 
b[20124] == 20124 && 
b[20125] == 20125 && 
b[20126] == 20126 && 
b[20127] == 20127 && 
b[20128] == 20128 && 
b[20129] == 20129 && 
b[20130] == 20130 && 
b[20131] == 20131 && 
b[20132] == 20132 && 
b[20133] == 20133 && 
b[20134] == 20134 && 
b[20135] == 20135 && 
b[20136] == 20136 && 
b[20137] == 20137 && 
b[20138] == 20138 && 
b[20139] == 20139 && 
b[20140] == 20140 && 
b[20141] == 20141 && 
b[20142] == 20142 && 
b[20143] == 20143 && 
b[20144] == 20144 && 
b[20145] == 20145 && 
b[20146] == 20146 && 
b[20147] == 20147 && 
b[20148] == 20148 && 
b[20149] == 20149 && 
b[20150] == 20150 && 
b[20151] == 20151 && 
b[20152] == 20152 && 
b[20153] == 20153 && 
b[20154] == 20154 && 
b[20155] == 20155 && 
b[20156] == 20156 && 
b[20157] == 20157 && 
b[20158] == 20158 && 
b[20159] == 20159 && 
b[20160] == 20160 && 
b[20161] == 20161 && 
b[20162] == 20162 && 
b[20163] == 20163 && 
b[20164] == 20164 && 
b[20165] == 20165 && 
b[20166] == 20166 && 
b[20167] == 20167 && 
b[20168] == 20168 && 
b[20169] == 20169 && 
b[20170] == 20170 && 
b[20171] == 20171 && 
b[20172] == 20172 && 
b[20173] == 20173 && 
b[20174] == 20174 && 
b[20175] == 20175 && 
b[20176] == 20176 && 
b[20177] == 20177 && 
b[20178] == 20178 && 
b[20179] == 20179 && 
b[20180] == 20180 && 
b[20181] == 20181 && 
b[20182] == 20182 && 
b[20183] == 20183 && 
b[20184] == 20184 && 
b[20185] == 20185 && 
b[20186] == 20186 && 
b[20187] == 20187 && 
b[20188] == 20188 && 
b[20189] == 20189 && 
b[20190] == 20190 && 
b[20191] == 20191 && 
b[20192] == 20192 && 
b[20193] == 20193 && 
b[20194] == 20194 && 
b[20195] == 20195 && 
b[20196] == 20196 && 
b[20197] == 20197 && 
b[20198] == 20198 && 
b[20199] == 20199 && 
b[20200] == 20200 && 
b[20201] == 20201 && 
b[20202] == 20202 && 
b[20203] == 20203 && 
b[20204] == 20204 && 
b[20205] == 20205 && 
b[20206] == 20206 && 
b[20207] == 20207 && 
b[20208] == 20208 && 
b[20209] == 20209 && 
b[20210] == 20210 && 
b[20211] == 20211 && 
b[20212] == 20212 && 
b[20213] == 20213 && 
b[20214] == 20214 && 
b[20215] == 20215 && 
b[20216] == 20216 && 
b[20217] == 20217 && 
b[20218] == 20218 && 
b[20219] == 20219 && 
b[20220] == 20220 && 
b[20221] == 20221 && 
b[20222] == 20222 && 
b[20223] == 20223 && 
b[20224] == 20224 && 
b[20225] == 20225 && 
b[20226] == 20226 && 
b[20227] == 20227 && 
b[20228] == 20228 && 
b[20229] == 20229 && 
b[20230] == 20230 && 
b[20231] == 20231 && 
b[20232] == 20232 && 
b[20233] == 20233 && 
b[20234] == 20234 && 
b[20235] == 20235 && 
b[20236] == 20236 && 
b[20237] == 20237 && 
b[20238] == 20238 && 
b[20239] == 20239 && 
b[20240] == 20240 && 
b[20241] == 20241 && 
b[20242] == 20242 && 
b[20243] == 20243 && 
b[20244] == 20244 && 
b[20245] == 20245 && 
b[20246] == 20246 && 
b[20247] == 20247 && 
b[20248] == 20248 && 
b[20249] == 20249 && 
b[20250] == 20250 && 
b[20251] == 20251 && 
b[20252] == 20252 && 
b[20253] == 20253 && 
b[20254] == 20254 && 
b[20255] == 20255 && 
b[20256] == 20256 && 
b[20257] == 20257 && 
b[20258] == 20258 && 
b[20259] == 20259 && 
b[20260] == 20260 && 
b[20261] == 20261 && 
b[20262] == 20262 && 
b[20263] == 20263 && 
b[20264] == 20264 && 
b[20265] == 20265 && 
b[20266] == 20266 && 
b[20267] == 20267 && 
b[20268] == 20268 && 
b[20269] == 20269 && 
b[20270] == 20270 && 
b[20271] == 20271 && 
b[20272] == 20272 && 
b[20273] == 20273 && 
b[20274] == 20274 && 
b[20275] == 20275 && 
b[20276] == 20276 && 
b[20277] == 20277 && 
b[20278] == 20278 && 
b[20279] == 20279 && 
b[20280] == 20280 && 
b[20281] == 20281 && 
b[20282] == 20282 && 
b[20283] == 20283 && 
b[20284] == 20284 && 
b[20285] == 20285 && 
b[20286] == 20286 && 
b[20287] == 20287 && 
b[20288] == 20288 && 
b[20289] == 20289 && 
b[20290] == 20290 && 
b[20291] == 20291 && 
b[20292] == 20292 && 
b[20293] == 20293 && 
b[20294] == 20294 && 
b[20295] == 20295 && 
b[20296] == 20296 && 
b[20297] == 20297 && 
b[20298] == 20298 && 
b[20299] == 20299 && 
b[20300] == 20300 && 
b[20301] == 20301 && 
b[20302] == 20302 && 
b[20303] == 20303 && 
b[20304] == 20304 && 
b[20305] == 20305 && 
b[20306] == 20306 && 
b[20307] == 20307 && 
b[20308] == 20308 && 
b[20309] == 20309 && 
b[20310] == 20310 && 
b[20311] == 20311 && 
b[20312] == 20312 && 
b[20313] == 20313 && 
b[20314] == 20314 && 
b[20315] == 20315 && 
b[20316] == 20316 && 
b[20317] == 20317 && 
b[20318] == 20318 && 
b[20319] == 20319 && 
b[20320] == 20320 && 
b[20321] == 20321 && 
b[20322] == 20322 && 
b[20323] == 20323 && 
b[20324] == 20324 && 
b[20325] == 20325 && 
b[20326] == 20326 && 
b[20327] == 20327 && 
b[20328] == 20328 && 
b[20329] == 20329 && 
b[20330] == 20330 && 
b[20331] == 20331 && 
b[20332] == 20332 && 
b[20333] == 20333 && 
b[20334] == 20334 && 
b[20335] == 20335 && 
b[20336] == 20336 && 
b[20337] == 20337 && 
b[20338] == 20338 && 
b[20339] == 20339 && 
b[20340] == 20340 && 
b[20341] == 20341 && 
b[20342] == 20342 && 
b[20343] == 20343 && 
b[20344] == 20344 && 
b[20345] == 20345 && 
b[20346] == 20346 && 
b[20347] == 20347 && 
b[20348] == 20348 && 
b[20349] == 20349 && 
b[20350] == 20350 && 
b[20351] == 20351 && 
b[20352] == 20352 && 
b[20353] == 20353 && 
b[20354] == 20354 && 
b[20355] == 20355 && 
b[20356] == 20356 && 
b[20357] == 20357 && 
b[20358] == 20358 && 
b[20359] == 20359 && 
b[20360] == 20360 && 
b[20361] == 20361 && 
b[20362] == 20362 && 
b[20363] == 20363 && 
b[20364] == 20364 && 
b[20365] == 20365 && 
b[20366] == 20366 && 
b[20367] == 20367 && 
b[20368] == 20368 && 
b[20369] == 20369 && 
b[20370] == 20370 && 
b[20371] == 20371 && 
b[20372] == 20372 && 
b[20373] == 20373 && 
b[20374] == 20374 && 
b[20375] == 20375 && 
b[20376] == 20376 && 
b[20377] == 20377 && 
b[20378] == 20378 && 
b[20379] == 20379 && 
b[20380] == 20380 && 
b[20381] == 20381 && 
b[20382] == 20382 && 
b[20383] == 20383 && 
b[20384] == 20384 && 
b[20385] == 20385 && 
b[20386] == 20386 && 
b[20387] == 20387 && 
b[20388] == 20388 && 
b[20389] == 20389 && 
b[20390] == 20390 && 
b[20391] == 20391 && 
b[20392] == 20392 && 
b[20393] == 20393 && 
b[20394] == 20394 && 
b[20395] == 20395 && 
b[20396] == 20396 && 
b[20397] == 20397 && 
b[20398] == 20398 && 
b[20399] == 20399 && 
b[20400] == 20400 && 
b[20401] == 20401 && 
b[20402] == 20402 && 
b[20403] == 20403 && 
b[20404] == 20404 && 
b[20405] == 20405 && 
b[20406] == 20406 && 
b[20407] == 20407 && 
b[20408] == 20408 && 
b[20409] == 20409 && 
b[20410] == 20410 && 
b[20411] == 20411 && 
b[20412] == 20412 && 
b[20413] == 20413 && 
b[20414] == 20414 && 
b[20415] == 20415 && 
b[20416] == 20416 && 
b[20417] == 20417 && 
b[20418] == 20418 && 
b[20419] == 20419 && 
b[20420] == 20420 && 
b[20421] == 20421 && 
b[20422] == 20422 && 
b[20423] == 20423 && 
b[20424] == 20424 && 
b[20425] == 20425 && 
b[20426] == 20426 && 
b[20427] == 20427 && 
b[20428] == 20428 && 
b[20429] == 20429 && 
b[20430] == 20430 && 
b[20431] == 20431 && 
b[20432] == 20432 && 
b[20433] == 20433 && 
b[20434] == 20434 && 
b[20435] == 20435 && 
b[20436] == 20436 && 
b[20437] == 20437 && 
b[20438] == 20438 && 
b[20439] == 20439 && 
b[20440] == 20440 && 
b[20441] == 20441 && 
b[20442] == 20442 && 
b[20443] == 20443 && 
b[20444] == 20444 && 
b[20445] == 20445 && 
b[20446] == 20446 && 
b[20447] == 20447 && 
b[20448] == 20448 && 
b[20449] == 20449 && 
b[20450] == 20450 && 
b[20451] == 20451 && 
b[20452] == 20452 && 
b[20453] == 20453 && 
b[20454] == 20454 && 
b[20455] == 20455 && 
b[20456] == 20456 && 
b[20457] == 20457 && 
b[20458] == 20458 && 
b[20459] == 20459 && 
b[20460] == 20460 && 
b[20461] == 20461 && 
b[20462] == 20462 && 
b[20463] == 20463 && 
b[20464] == 20464 && 
b[20465] == 20465 && 
b[20466] == 20466 && 
b[20467] == 20467 && 
b[20468] == 20468 && 
b[20469] == 20469 && 
b[20470] == 20470 && 
b[20471] == 20471 && 
b[20472] == 20472 && 
b[20473] == 20473 && 
b[20474] == 20474 && 
b[20475] == 20475 && 
b[20476] == 20476 && 
b[20477] == 20477 && 
b[20478] == 20478 && 
b[20479] == 20479 && 
b[20480] == 20480 && 
b[20481] == 20481 && 
b[20482] == 20482 && 
b[20483] == 20483 && 
b[20484] == 20484 && 
b[20485] == 20485 && 
b[20486] == 20486 && 
b[20487] == 20487 && 
b[20488] == 20488 && 
b[20489] == 20489 && 
b[20490] == 20490 && 
b[20491] == 20491 && 
b[20492] == 20492 && 
b[20493] == 20493 && 
b[20494] == 20494 && 
b[20495] == 20495 && 
b[20496] == 20496 && 
b[20497] == 20497 && 
b[20498] == 20498 && 
b[20499] == 20499 && 
b[20500] == 20500 && 
b[20501] == 20501 && 
b[20502] == 20502 && 
b[20503] == 20503 && 
b[20504] == 20504 && 
b[20505] == 20505 && 
b[20506] == 20506 && 
b[20507] == 20507 && 
b[20508] == 20508 && 
b[20509] == 20509 && 
b[20510] == 20510 && 
b[20511] == 20511 && 
b[20512] == 20512 && 
b[20513] == 20513 && 
b[20514] == 20514 && 
b[20515] == 20515 && 
b[20516] == 20516 && 
b[20517] == 20517 && 
b[20518] == 20518 && 
b[20519] == 20519 && 
b[20520] == 20520 && 
b[20521] == 20521 && 
b[20522] == 20522 && 
b[20523] == 20523 && 
b[20524] == 20524 && 
b[20525] == 20525 && 
b[20526] == 20526 && 
b[20527] == 20527 && 
b[20528] == 20528 && 
b[20529] == 20529 && 
b[20530] == 20530 && 
b[20531] == 20531 && 
b[20532] == 20532 && 
b[20533] == 20533 && 
b[20534] == 20534 && 
b[20535] == 20535 && 
b[20536] == 20536 && 
b[20537] == 20537 && 
b[20538] == 20538 && 
b[20539] == 20539 && 
b[20540] == 20540 && 
b[20541] == 20541 && 
b[20542] == 20542 && 
b[20543] == 20543 && 
b[20544] == 20544 && 
b[20545] == 20545 && 
b[20546] == 20546 && 
b[20547] == 20547 && 
b[20548] == 20548 && 
b[20549] == 20549 && 
b[20550] == 20550 && 
b[20551] == 20551 && 
b[20552] == 20552 && 
b[20553] == 20553 && 
b[20554] == 20554 && 
b[20555] == 20555 && 
b[20556] == 20556 && 
b[20557] == 20557 && 
b[20558] == 20558 && 
b[20559] == 20559 && 
b[20560] == 20560 && 
b[20561] == 20561 && 
b[20562] == 20562 && 
b[20563] == 20563 && 
b[20564] == 20564 && 
b[20565] == 20565 && 
b[20566] == 20566 && 
b[20567] == 20567 && 
b[20568] == 20568 && 
b[20569] == 20569 && 
b[20570] == 20570 && 
b[20571] == 20571 && 
b[20572] == 20572 && 
b[20573] == 20573 && 
b[20574] == 20574 && 
b[20575] == 20575 && 
b[20576] == 20576 && 
b[20577] == 20577 && 
b[20578] == 20578 && 
b[20579] == 20579 && 
b[20580] == 20580 && 
b[20581] == 20581 && 
b[20582] == 20582 && 
b[20583] == 20583 && 
b[20584] == 20584 && 
b[20585] == 20585 && 
b[20586] == 20586 && 
b[20587] == 20587 && 
b[20588] == 20588 && 
b[20589] == 20589 && 
b[20590] == 20590 && 
b[20591] == 20591 && 
b[20592] == 20592 && 
b[20593] == 20593 && 
b[20594] == 20594 && 
b[20595] == 20595 && 
b[20596] == 20596 && 
b[20597] == 20597 && 
b[20598] == 20598 && 
b[20599] == 20599 && 
b[20600] == 20600 && 
b[20601] == 20601 && 
b[20602] == 20602 && 
b[20603] == 20603 && 
b[20604] == 20604 && 
b[20605] == 20605 && 
b[20606] == 20606 && 
b[20607] == 20607 && 
b[20608] == 20608 && 
b[20609] == 20609 && 
b[20610] == 20610 && 
b[20611] == 20611 && 
b[20612] == 20612 && 
b[20613] == 20613 && 
b[20614] == 20614 && 
b[20615] == 20615 && 
b[20616] == 20616 && 
b[20617] == 20617 && 
b[20618] == 20618 && 
b[20619] == 20619 && 
b[20620] == 20620 && 
b[20621] == 20621 && 
b[20622] == 20622 && 
b[20623] == 20623 && 
b[20624] == 20624 && 
b[20625] == 20625 && 
b[20626] == 20626 && 
b[20627] == 20627 && 
b[20628] == 20628 && 
b[20629] == 20629 && 
b[20630] == 20630 && 
b[20631] == 20631 && 
b[20632] == 20632 && 
b[20633] == 20633 && 
b[20634] == 20634 && 
b[20635] == 20635 && 
b[20636] == 20636 && 
b[20637] == 20637 && 
b[20638] == 20638 && 
b[20639] == 20639 && 
b[20640] == 20640 && 
b[20641] == 20641 && 
b[20642] == 20642 && 
b[20643] == 20643 && 
b[20644] == 20644 && 
b[20645] == 20645 && 
b[20646] == 20646 && 
b[20647] == 20647 && 
b[20648] == 20648 && 
b[20649] == 20649 && 
b[20650] == 20650 && 
b[20651] == 20651 && 
b[20652] == 20652 && 
b[20653] == 20653 && 
b[20654] == 20654 && 
b[20655] == 20655 && 
b[20656] == 20656 && 
b[20657] == 20657 && 
b[20658] == 20658 && 
b[20659] == 20659 && 
b[20660] == 20660 && 
b[20661] == 20661 && 
b[20662] == 20662 && 
b[20663] == 20663 && 
b[20664] == 20664 && 
b[20665] == 20665 && 
b[20666] == 20666 && 
b[20667] == 20667 && 
b[20668] == 20668 && 
b[20669] == 20669 && 
b[20670] == 20670 && 
b[20671] == 20671 && 
b[20672] == 20672 && 
b[20673] == 20673 && 
b[20674] == 20674 && 
b[20675] == 20675 && 
b[20676] == 20676 && 
b[20677] == 20677 && 
b[20678] == 20678 && 
b[20679] == 20679 && 
b[20680] == 20680 && 
b[20681] == 20681 && 
b[20682] == 20682 && 
b[20683] == 20683 && 
b[20684] == 20684 && 
b[20685] == 20685 && 
b[20686] == 20686 && 
b[20687] == 20687 && 
b[20688] == 20688 && 
b[20689] == 20689 && 
b[20690] == 20690 && 
b[20691] == 20691 && 
b[20692] == 20692 && 
b[20693] == 20693 && 
b[20694] == 20694 && 
b[20695] == 20695 && 
b[20696] == 20696 && 
b[20697] == 20697 && 
b[20698] == 20698 && 
b[20699] == 20699 && 
b[20700] == 20700 && 
b[20701] == 20701 && 
b[20702] == 20702 && 
b[20703] == 20703 && 
b[20704] == 20704 && 
b[20705] == 20705 && 
b[20706] == 20706 && 
b[20707] == 20707 && 
b[20708] == 20708 && 
b[20709] == 20709 && 
b[20710] == 20710 && 
b[20711] == 20711 && 
b[20712] == 20712 && 
b[20713] == 20713 && 
b[20714] == 20714 && 
b[20715] == 20715 && 
b[20716] == 20716 && 
b[20717] == 20717 && 
b[20718] == 20718 && 
b[20719] == 20719 && 
b[20720] == 20720 && 
b[20721] == 20721 && 
b[20722] == 20722 && 
b[20723] == 20723 && 
b[20724] == 20724 && 
b[20725] == 20725 && 
b[20726] == 20726 && 
b[20727] == 20727 && 
b[20728] == 20728 && 
b[20729] == 20729 && 
b[20730] == 20730 && 
b[20731] == 20731 && 
b[20732] == 20732 && 
b[20733] == 20733 && 
b[20734] == 20734 && 
b[20735] == 20735 && 
b[20736] == 20736 && 
b[20737] == 20737 && 
b[20738] == 20738 && 
b[20739] == 20739 && 
b[20740] == 20740 && 
b[20741] == 20741 && 
b[20742] == 20742 && 
b[20743] == 20743 && 
b[20744] == 20744 && 
b[20745] == 20745 && 
b[20746] == 20746 && 
b[20747] == 20747 && 
b[20748] == 20748 && 
b[20749] == 20749 && 
b[20750] == 20750 && 
b[20751] == 20751 && 
b[20752] == 20752 && 
b[20753] == 20753 && 
b[20754] == 20754 && 
b[20755] == 20755 && 
b[20756] == 20756 && 
b[20757] == 20757 && 
b[20758] == 20758 && 
b[20759] == 20759 && 
b[20760] == 20760 && 
b[20761] == 20761 && 
b[20762] == 20762 && 
b[20763] == 20763 && 
b[20764] == 20764 && 
b[20765] == 20765 && 
b[20766] == 20766 && 
b[20767] == 20767 && 
b[20768] == 20768 && 
b[20769] == 20769 && 
b[20770] == 20770 && 
b[20771] == 20771 && 
b[20772] == 20772 && 
b[20773] == 20773 && 
b[20774] == 20774 && 
b[20775] == 20775 && 
b[20776] == 20776 && 
b[20777] == 20777 && 
b[20778] == 20778 && 
b[20779] == 20779 && 
b[20780] == 20780 && 
b[20781] == 20781 && 
b[20782] == 20782 && 
b[20783] == 20783 && 
b[20784] == 20784 && 
b[20785] == 20785 && 
b[20786] == 20786 && 
b[20787] == 20787 && 
b[20788] == 20788 && 
b[20789] == 20789 && 
b[20790] == 20790 && 
b[20791] == 20791 && 
b[20792] == 20792 && 
b[20793] == 20793 && 
b[20794] == 20794 && 
b[20795] == 20795 && 
b[20796] == 20796 && 
b[20797] == 20797 && 
b[20798] == 20798 && 
b[20799] == 20799 && 
b[20800] == 20800 && 
b[20801] == 20801 && 
b[20802] == 20802 && 
b[20803] == 20803 && 
b[20804] == 20804 && 
b[20805] == 20805 && 
b[20806] == 20806 && 
b[20807] == 20807 && 
b[20808] == 20808 && 
b[20809] == 20809 && 
b[20810] == 20810 && 
b[20811] == 20811 && 
b[20812] == 20812 && 
b[20813] == 20813 && 
b[20814] == 20814 && 
b[20815] == 20815 && 
b[20816] == 20816 && 
b[20817] == 20817 && 
b[20818] == 20818 && 
b[20819] == 20819 && 
b[20820] == 20820 && 
b[20821] == 20821 && 
b[20822] == 20822 && 
b[20823] == 20823 && 
b[20824] == 20824 && 
b[20825] == 20825 && 
b[20826] == 20826 && 
b[20827] == 20827 && 
b[20828] == 20828 && 
b[20829] == 20829 && 
b[20830] == 20830 && 
b[20831] == 20831 && 
b[20832] == 20832 && 
b[20833] == 20833 && 
b[20834] == 20834 && 
b[20835] == 20835 && 
b[20836] == 20836 && 
b[20837] == 20837 && 
b[20838] == 20838 && 
b[20839] == 20839 && 
b[20840] == 20840 && 
b[20841] == 20841 && 
b[20842] == 20842 && 
b[20843] == 20843 && 
b[20844] == 20844 && 
b[20845] == 20845 && 
b[20846] == 20846 && 
b[20847] == 20847 && 
b[20848] == 20848 && 
b[20849] == 20849 && 
b[20850] == 20850 && 
b[20851] == 20851 && 
b[20852] == 20852 && 
b[20853] == 20853 && 
b[20854] == 20854 && 
b[20855] == 20855 && 
b[20856] == 20856 && 
b[20857] == 20857 && 
b[20858] == 20858 && 
b[20859] == 20859 && 
b[20860] == 20860 && 
b[20861] == 20861 && 
b[20862] == 20862 && 
b[20863] == 20863 && 
b[20864] == 20864 && 
b[20865] == 20865 && 
b[20866] == 20866 && 
b[20867] == 20867 && 
b[20868] == 20868 && 
b[20869] == 20869 && 
b[20870] == 20870 && 
b[20871] == 20871 && 
b[20872] == 20872 && 
b[20873] == 20873 && 
b[20874] == 20874 && 
b[20875] == 20875 && 
b[20876] == 20876 && 
b[20877] == 20877 && 
b[20878] == 20878 && 
b[20879] == 20879 && 
b[20880] == 20880 && 
b[20881] == 20881 && 
b[20882] == 20882 && 
b[20883] == 20883 && 
b[20884] == 20884 && 
b[20885] == 20885 && 
b[20886] == 20886 && 
b[20887] == 20887 && 
b[20888] == 20888 && 
b[20889] == 20889 && 
b[20890] == 20890 && 
b[20891] == 20891 && 
b[20892] == 20892 && 
b[20893] == 20893 && 
b[20894] == 20894 && 
b[20895] == 20895 && 
b[20896] == 20896 && 
b[20897] == 20897 && 
b[20898] == 20898 && 
b[20899] == 20899 && 
b[20900] == 20900 && 
b[20901] == 20901 && 
b[20902] == 20902 && 
b[20903] == 20903 && 
b[20904] == 20904 && 
b[20905] == 20905 && 
b[20906] == 20906 && 
b[20907] == 20907 && 
b[20908] == 20908 && 
b[20909] == 20909 && 
b[20910] == 20910 && 
b[20911] == 20911 && 
b[20912] == 20912 && 
b[20913] == 20913 && 
b[20914] == 20914 && 
b[20915] == 20915 && 
b[20916] == 20916 && 
b[20917] == 20917 && 
b[20918] == 20918 && 
b[20919] == 20919 && 
b[20920] == 20920 && 
b[20921] == 20921 && 
b[20922] == 20922 && 
b[20923] == 20923 && 
b[20924] == 20924 && 
b[20925] == 20925 && 
b[20926] == 20926 && 
b[20927] == 20927 && 
b[20928] == 20928 && 
b[20929] == 20929 && 
b[20930] == 20930 && 
b[20931] == 20931 && 
b[20932] == 20932 && 
b[20933] == 20933 && 
b[20934] == 20934 && 
b[20935] == 20935 && 
b[20936] == 20936 && 
b[20937] == 20937 && 
b[20938] == 20938 && 
b[20939] == 20939 && 
b[20940] == 20940 && 
b[20941] == 20941 && 
b[20942] == 20942 && 
b[20943] == 20943 && 
b[20944] == 20944 && 
b[20945] == 20945 && 
b[20946] == 20946 && 
b[20947] == 20947 && 
b[20948] == 20948 && 
b[20949] == 20949 && 
b[20950] == 20950 && 
b[20951] == 20951 && 
b[20952] == 20952 && 
b[20953] == 20953 && 
b[20954] == 20954 && 
b[20955] == 20955 && 
b[20956] == 20956 && 
b[20957] == 20957 && 
b[20958] == 20958 && 
b[20959] == 20959 && 
b[20960] == 20960 && 
b[20961] == 20961 && 
b[20962] == 20962 && 
b[20963] == 20963 && 
b[20964] == 20964 && 
b[20965] == 20965 && 
b[20966] == 20966 && 
b[20967] == 20967 && 
b[20968] == 20968 && 
b[20969] == 20969 && 
b[20970] == 20970 && 
b[20971] == 20971 && 
b[20972] == 20972 && 
b[20973] == 20973 && 
b[20974] == 20974 && 
b[20975] == 20975 && 
b[20976] == 20976 && 
b[20977] == 20977 && 
b[20978] == 20978 && 
b[20979] == 20979 && 
b[20980] == 20980 && 
b[20981] == 20981 && 
b[20982] == 20982 && 
b[20983] == 20983 && 
b[20984] == 20984 && 
b[20985] == 20985 && 
b[20986] == 20986 && 
b[20987] == 20987 && 
b[20988] == 20988 && 
b[20989] == 20989 && 
b[20990] == 20990 && 
b[20991] == 20991 && 
b[20992] == 20992 && 
b[20993] == 20993 && 
b[20994] == 20994 && 
b[20995] == 20995 && 
b[20996] == 20996 && 
b[20997] == 20997 && 
b[20998] == 20998 && 
b[20999] == 20999 && 
b[21000] == 21000 && 
b[21001] == 21001 && 
b[21002] == 21002 && 
b[21003] == 21003 && 
b[21004] == 21004 && 
b[21005] == 21005 && 
b[21006] == 21006 && 
b[21007] == 21007 && 
b[21008] == 21008 && 
b[21009] == 21009 && 
b[21010] == 21010 && 
b[21011] == 21011 && 
b[21012] == 21012 && 
b[21013] == 21013 && 
b[21014] == 21014 && 
b[21015] == 21015 && 
b[21016] == 21016 && 
b[21017] == 21017 && 
b[21018] == 21018 && 
b[21019] == 21019 && 
b[21020] == 21020 && 
b[21021] == 21021 && 
b[21022] == 21022 && 
b[21023] == 21023 && 
b[21024] == 21024 && 
b[21025] == 21025 && 
b[21026] == 21026 && 
b[21027] == 21027 && 
b[21028] == 21028 && 
b[21029] == 21029 && 
b[21030] == 21030 && 
b[21031] == 21031 && 
b[21032] == 21032 && 
b[21033] == 21033 && 
b[21034] == 21034 && 
b[21035] == 21035 && 
b[21036] == 21036 && 
b[21037] == 21037 && 
b[21038] == 21038 && 
b[21039] == 21039 && 
b[21040] == 21040 && 
b[21041] == 21041 && 
b[21042] == 21042 && 
b[21043] == 21043 && 
b[21044] == 21044 && 
b[21045] == 21045 && 
b[21046] == 21046 && 
b[21047] == 21047 && 
b[21048] == 21048 && 
b[21049] == 21049 && 
b[21050] == 21050 && 
b[21051] == 21051 && 
b[21052] == 21052 && 
b[21053] == 21053 && 
b[21054] == 21054 && 
b[21055] == 21055 && 
b[21056] == 21056 && 
b[21057] == 21057 && 
b[21058] == 21058 && 
b[21059] == 21059 && 
b[21060] == 21060 && 
b[21061] == 21061 && 
b[21062] == 21062 && 
b[21063] == 21063 && 
b[21064] == 21064 && 
b[21065] == 21065 && 
b[21066] == 21066 && 
b[21067] == 21067 && 
b[21068] == 21068 && 
b[21069] == 21069 && 
b[21070] == 21070 && 
b[21071] == 21071 && 
b[21072] == 21072 && 
b[21073] == 21073 && 
b[21074] == 21074 && 
b[21075] == 21075 && 
b[21076] == 21076 && 
b[21077] == 21077 && 
b[21078] == 21078 && 
b[21079] == 21079 && 
b[21080] == 21080 && 
b[21081] == 21081 && 
b[21082] == 21082 && 
b[21083] == 21083 && 
b[21084] == 21084 && 
b[21085] == 21085 && 
b[21086] == 21086 && 
b[21087] == 21087 && 
b[21088] == 21088 && 
b[21089] == 21089 && 
b[21090] == 21090 && 
b[21091] == 21091 && 
b[21092] == 21092 && 
b[21093] == 21093 && 
b[21094] == 21094 && 
b[21095] == 21095 && 
b[21096] == 21096 && 
b[21097] == 21097 && 
b[21098] == 21098 && 
b[21099] == 21099 && 
b[21100] == 21100 && 
b[21101] == 21101 && 
b[21102] == 21102 && 
b[21103] == 21103 && 
b[21104] == 21104 && 
b[21105] == 21105 && 
b[21106] == 21106 && 
b[21107] == 21107 && 
b[21108] == 21108 && 
b[21109] == 21109 && 
b[21110] == 21110 && 
b[21111] == 21111 && 
b[21112] == 21112 && 
b[21113] == 21113 && 
b[21114] == 21114 && 
b[21115] == 21115 && 
b[21116] == 21116 && 
b[21117] == 21117 && 
b[21118] == 21118 && 
b[21119] == 21119 && 
b[21120] == 21120 && 
b[21121] == 21121 && 
b[21122] == 21122 && 
b[21123] == 21123 && 
b[21124] == 21124 && 
b[21125] == 21125 && 
b[21126] == 21126 && 
b[21127] == 21127 && 
b[21128] == 21128 && 
b[21129] == 21129 && 
b[21130] == 21130 && 
b[21131] == 21131 && 
b[21132] == 21132 && 
b[21133] == 21133 && 
b[21134] == 21134 && 
b[21135] == 21135 && 
b[21136] == 21136 && 
b[21137] == 21137 && 
b[21138] == 21138 && 
b[21139] == 21139 && 
b[21140] == 21140 && 
b[21141] == 21141 && 
b[21142] == 21142 && 
b[21143] == 21143 && 
b[21144] == 21144 && 
b[21145] == 21145 && 
b[21146] == 21146 && 
b[21147] == 21147 && 
b[21148] == 21148 && 
b[21149] == 21149 && 
b[21150] == 21150 && 
b[21151] == 21151 && 
b[21152] == 21152 && 
b[21153] == 21153 && 
b[21154] == 21154 && 
b[21155] == 21155 && 
b[21156] == 21156 && 
b[21157] == 21157 && 
b[21158] == 21158 && 
b[21159] == 21159 && 
b[21160] == 21160 && 
b[21161] == 21161 && 
b[21162] == 21162 && 
b[21163] == 21163 && 
b[21164] == 21164 && 
b[21165] == 21165 && 
b[21166] == 21166 && 
b[21167] == 21167 && 
b[21168] == 21168 && 
b[21169] == 21169 && 
b[21170] == 21170 && 
b[21171] == 21171 && 
b[21172] == 21172 && 
b[21173] == 21173 && 
b[21174] == 21174 && 
b[21175] == 21175 && 
b[21176] == 21176 && 
b[21177] == 21177 && 
b[21178] == 21178 && 
b[21179] == 21179 && 
b[21180] == 21180 && 
b[21181] == 21181 && 
b[21182] == 21182 && 
b[21183] == 21183 && 
b[21184] == 21184 && 
b[21185] == 21185 && 
b[21186] == 21186 && 
b[21187] == 21187 && 
b[21188] == 21188 && 
b[21189] == 21189 && 
b[21190] == 21190 && 
b[21191] == 21191 && 
b[21192] == 21192 && 
b[21193] == 21193 && 
b[21194] == 21194 && 
b[21195] == 21195 && 
b[21196] == 21196 && 
b[21197] == 21197 && 
b[21198] == 21198 && 
b[21199] == 21199 && 
b[21200] == 21200 && 
b[21201] == 21201 && 
b[21202] == 21202 && 
b[21203] == 21203 && 
b[21204] == 21204 && 
b[21205] == 21205 && 
b[21206] == 21206 && 
b[21207] == 21207 && 
b[21208] == 21208 && 
b[21209] == 21209 && 
b[21210] == 21210 && 
b[21211] == 21211 && 
b[21212] == 21212 && 
b[21213] == 21213 && 
b[21214] == 21214 && 
b[21215] == 21215 && 
b[21216] == 21216 && 
b[21217] == 21217 && 
b[21218] == 21218 && 
b[21219] == 21219 && 
b[21220] == 21220 && 
b[21221] == 21221 && 
b[21222] == 21222 && 
b[21223] == 21223 && 
b[21224] == 21224 && 
b[21225] == 21225 && 
b[21226] == 21226 && 
b[21227] == 21227 && 
b[21228] == 21228 && 
b[21229] == 21229 && 
b[21230] == 21230 && 
b[21231] == 21231 && 
b[21232] == 21232 && 
b[21233] == 21233 && 
b[21234] == 21234 && 
b[21235] == 21235 && 
b[21236] == 21236 && 
b[21237] == 21237 && 
b[21238] == 21238 && 
b[21239] == 21239 && 
b[21240] == 21240 && 
b[21241] == 21241 && 
b[21242] == 21242 && 
b[21243] == 21243 && 
b[21244] == 21244 && 
b[21245] == 21245 && 
b[21246] == 21246 && 
b[21247] == 21247 && 
b[21248] == 21248 && 
b[21249] == 21249 && 
b[21250] == 21250 && 
b[21251] == 21251 && 
b[21252] == 21252 && 
b[21253] == 21253 && 
b[21254] == 21254 && 
b[21255] == 21255 && 
b[21256] == 21256 && 
b[21257] == 21257 && 
b[21258] == 21258 && 
b[21259] == 21259 && 
b[21260] == 21260 && 
b[21261] == 21261 && 
b[21262] == 21262 && 
b[21263] == 21263 && 
b[21264] == 21264 && 
b[21265] == 21265 && 
b[21266] == 21266 && 
b[21267] == 21267 && 
b[21268] == 21268 && 
b[21269] == 21269 && 
b[21270] == 21270 && 
b[21271] == 21271 && 
b[21272] == 21272 && 
b[21273] == 21273 && 
b[21274] == 21274 && 
b[21275] == 21275 && 
b[21276] == 21276 && 
b[21277] == 21277 && 
b[21278] == 21278 && 
b[21279] == 21279 && 
b[21280] == 21280 && 
b[21281] == 21281 && 
b[21282] == 21282 && 
b[21283] == 21283 && 
b[21284] == 21284 && 
b[21285] == 21285 && 
b[21286] == 21286 && 
b[21287] == 21287 && 
b[21288] == 21288 && 
b[21289] == 21289 && 
b[21290] == 21290 && 
b[21291] == 21291 && 
b[21292] == 21292 && 
b[21293] == 21293 && 
b[21294] == 21294 && 
b[21295] == 21295 && 
b[21296] == 21296 && 
b[21297] == 21297 && 
b[21298] == 21298 && 
b[21299] == 21299 && 
b[21300] == 21300 && 
b[21301] == 21301 && 
b[21302] == 21302 && 
b[21303] == 21303 && 
b[21304] == 21304 && 
b[21305] == 21305 && 
b[21306] == 21306 && 
b[21307] == 21307 && 
b[21308] == 21308 && 
b[21309] == 21309 && 
b[21310] == 21310 && 
b[21311] == 21311 && 
b[21312] == 21312 && 
b[21313] == 21313 && 
b[21314] == 21314 && 
b[21315] == 21315 && 
b[21316] == 21316 && 
b[21317] == 21317 && 
b[21318] == 21318 && 
b[21319] == 21319 && 
b[21320] == 21320 && 
b[21321] == 21321 && 
b[21322] == 21322 && 
b[21323] == 21323 && 
b[21324] == 21324 && 
b[21325] == 21325 && 
b[21326] == 21326 && 
b[21327] == 21327 && 
b[21328] == 21328 && 
b[21329] == 21329 && 
b[21330] == 21330 && 
b[21331] == 21331 && 
b[21332] == 21332 && 
b[21333] == 21333 && 
b[21334] == 21334 && 
b[21335] == 21335 && 
b[21336] == 21336 && 
b[21337] == 21337 && 
b[21338] == 21338 && 
b[21339] == 21339 && 
b[21340] == 21340 && 
b[21341] == 21341 && 
b[21342] == 21342 && 
b[21343] == 21343 && 
b[21344] == 21344 && 
b[21345] == 21345 && 
b[21346] == 21346 && 
b[21347] == 21347 && 
b[21348] == 21348 && 
b[21349] == 21349 && 
b[21350] == 21350 && 
b[21351] == 21351 && 
b[21352] == 21352 && 
b[21353] == 21353 && 
b[21354] == 21354 && 
b[21355] == 21355 && 
b[21356] == 21356 && 
b[21357] == 21357 && 
b[21358] == 21358 && 
b[21359] == 21359 && 
b[21360] == 21360 && 
b[21361] == 21361 && 
b[21362] == 21362 && 
b[21363] == 21363 && 
b[21364] == 21364 && 
b[21365] == 21365 && 
b[21366] == 21366 && 
b[21367] == 21367 && 
b[21368] == 21368 && 
b[21369] == 21369 && 
b[21370] == 21370 && 
b[21371] == 21371 && 
b[21372] == 21372 && 
b[21373] == 21373 && 
b[21374] == 21374 && 
b[21375] == 21375 && 
b[21376] == 21376 && 
b[21377] == 21377 && 
b[21378] == 21378 && 
b[21379] == 21379 && 
b[21380] == 21380 && 
b[21381] == 21381 && 
b[21382] == 21382 && 
b[21383] == 21383 && 
b[21384] == 21384 && 
b[21385] == 21385 && 
b[21386] == 21386 && 
b[21387] == 21387 && 
b[21388] == 21388 && 
b[21389] == 21389 && 
b[21390] == 21390 && 
b[21391] == 21391 && 
b[21392] == 21392 && 
b[21393] == 21393 && 
b[21394] == 21394 && 
b[21395] == 21395 && 
b[21396] == 21396 && 
b[21397] == 21397 && 
b[21398] == 21398 && 
b[21399] == 21399 && 
b[21400] == 21400 && 
b[21401] == 21401 && 
b[21402] == 21402 && 
b[21403] == 21403 && 
b[21404] == 21404 && 
b[21405] == 21405 && 
b[21406] == 21406 && 
b[21407] == 21407 && 
b[21408] == 21408 && 
b[21409] == 21409 && 
b[21410] == 21410 && 
b[21411] == 21411 && 
b[21412] == 21412 && 
b[21413] == 21413 && 
b[21414] == 21414 && 
b[21415] == 21415 && 
b[21416] == 21416 && 
b[21417] == 21417 && 
b[21418] == 21418 && 
b[21419] == 21419 && 
b[21420] == 21420 && 
b[21421] == 21421 && 
b[21422] == 21422 && 
b[21423] == 21423 && 
b[21424] == 21424 && 
b[21425] == 21425 && 
b[21426] == 21426 && 
b[21427] == 21427 && 
b[21428] == 21428 && 
b[21429] == 21429 && 
b[21430] == 21430 && 
b[21431] == 21431 && 
b[21432] == 21432 && 
b[21433] == 21433 && 
b[21434] == 21434 && 
b[21435] == 21435 && 
b[21436] == 21436 && 
b[21437] == 21437 && 
b[21438] == 21438 && 
b[21439] == 21439 && 
b[21440] == 21440 && 
b[21441] == 21441 && 
b[21442] == 21442 && 
b[21443] == 21443 && 
b[21444] == 21444 && 
b[21445] == 21445 && 
b[21446] == 21446 && 
b[21447] == 21447 && 
b[21448] == 21448 && 
b[21449] == 21449 && 
b[21450] == 21450 && 
b[21451] == 21451 && 
b[21452] == 21452 && 
b[21453] == 21453 && 
b[21454] == 21454 && 
b[21455] == 21455 && 
b[21456] == 21456 && 
b[21457] == 21457 && 
b[21458] == 21458 && 
b[21459] == 21459 && 
b[21460] == 21460 && 
b[21461] == 21461 && 
b[21462] == 21462 && 
b[21463] == 21463 && 
b[21464] == 21464 && 
b[21465] == 21465 && 
b[21466] == 21466 && 
b[21467] == 21467 && 
b[21468] == 21468 && 
b[21469] == 21469 && 
b[21470] == 21470 && 
b[21471] == 21471 && 
b[21472] == 21472 && 
b[21473] == 21473 && 
b[21474] == 21474 && 
b[21475] == 21475 && 
b[21476] == 21476 && 
b[21477] == 21477 && 
b[21478] == 21478 && 
b[21479] == 21479 && 
b[21480] == 21480 && 
b[21481] == 21481 && 
b[21482] == 21482 && 
b[21483] == 21483 && 
b[21484] == 21484 && 
b[21485] == 21485 && 
b[21486] == 21486 && 
b[21487] == 21487 && 
b[21488] == 21488 && 
b[21489] == 21489 && 
b[21490] == 21490 && 
b[21491] == 21491 && 
b[21492] == 21492 && 
b[21493] == 21493 && 
b[21494] == 21494 && 
b[21495] == 21495 && 
b[21496] == 21496 && 
b[21497] == 21497 && 
b[21498] == 21498 && 
b[21499] == 21499 && 
b[21500] == 21500 && 
b[21501] == 21501 && 
b[21502] == 21502 && 
b[21503] == 21503 && 
b[21504] == 21504 && 
b[21505] == 21505 && 
b[21506] == 21506 && 
b[21507] == 21507 && 
b[21508] == 21508 && 
b[21509] == 21509 && 
b[21510] == 21510 && 
b[21511] == 21511 && 
b[21512] == 21512 && 
b[21513] == 21513 && 
b[21514] == 21514 && 
b[21515] == 21515 && 
b[21516] == 21516 && 
b[21517] == 21517 && 
b[21518] == 21518 && 
b[21519] == 21519 && 
b[21520] == 21520 && 
b[21521] == 21521 && 
b[21522] == 21522 && 
b[21523] == 21523 && 
b[21524] == 21524 && 
b[21525] == 21525 && 
b[21526] == 21526 && 
b[21527] == 21527 && 
b[21528] == 21528 && 
b[21529] == 21529 && 
b[21530] == 21530 && 
b[21531] == 21531 && 
b[21532] == 21532 && 
b[21533] == 21533 && 
b[21534] == 21534 && 
b[21535] == 21535 && 
b[21536] == 21536 && 
b[21537] == 21537 && 
b[21538] == 21538 && 
b[21539] == 21539 && 
b[21540] == 21540 && 
b[21541] == 21541 && 
b[21542] == 21542 && 
b[21543] == 21543 && 
b[21544] == 21544 && 
b[21545] == 21545 && 
b[21546] == 21546 && 
b[21547] == 21547 && 
b[21548] == 21548 && 
b[21549] == 21549 && 
b[21550] == 21550 && 
b[21551] == 21551 && 
b[21552] == 21552 && 
b[21553] == 21553 && 
b[21554] == 21554 && 
b[21555] == 21555 && 
b[21556] == 21556 && 
b[21557] == 21557 && 
b[21558] == 21558 && 
b[21559] == 21559 && 
b[21560] == 21560 && 
b[21561] == 21561 && 
b[21562] == 21562 && 
b[21563] == 21563 && 
b[21564] == 21564 && 
b[21565] == 21565 && 
b[21566] == 21566 && 
b[21567] == 21567 && 
b[21568] == 21568 && 
b[21569] == 21569 && 
b[21570] == 21570 && 
b[21571] == 21571 && 
b[21572] == 21572 && 
b[21573] == 21573 && 
b[21574] == 21574 && 
b[21575] == 21575 && 
b[21576] == 21576 && 
b[21577] == 21577 && 
b[21578] == 21578 && 
b[21579] == 21579 && 
b[21580] == 21580 && 
b[21581] == 21581 && 
b[21582] == 21582 && 
b[21583] == 21583 && 
b[21584] == 21584 && 
b[21585] == 21585 && 
b[21586] == 21586 && 
b[21587] == 21587 && 
b[21588] == 21588 && 
b[21589] == 21589 && 
b[21590] == 21590 && 
b[21591] == 21591 && 
b[21592] == 21592 && 
b[21593] == 21593 && 
b[21594] == 21594 && 
b[21595] == 21595 && 
b[21596] == 21596 && 
b[21597] == 21597 && 
b[21598] == 21598 && 
b[21599] == 21599 && 
b[21600] == 21600 && 
b[21601] == 21601 && 
b[21602] == 21602 && 
b[21603] == 21603 && 
b[21604] == 21604 && 
b[21605] == 21605 && 
b[21606] == 21606 && 
b[21607] == 21607 && 
b[21608] == 21608 && 
b[21609] == 21609 && 
b[21610] == 21610 && 
b[21611] == 21611 && 
b[21612] == 21612 && 
b[21613] == 21613 && 
b[21614] == 21614 && 
b[21615] == 21615 && 
b[21616] == 21616 && 
b[21617] == 21617 && 
b[21618] == 21618 && 
b[21619] == 21619 && 
b[21620] == 21620 && 
b[21621] == 21621 && 
b[21622] == 21622 && 
b[21623] == 21623 && 
b[21624] == 21624 && 
b[21625] == 21625 && 
b[21626] == 21626 && 
b[21627] == 21627 && 
b[21628] == 21628 && 
b[21629] == 21629 && 
b[21630] == 21630 && 
b[21631] == 21631 && 
b[21632] == 21632 && 
b[21633] == 21633 && 
b[21634] == 21634 && 
b[21635] == 21635 && 
b[21636] == 21636 && 
b[21637] == 21637 && 
b[21638] == 21638 && 
b[21639] == 21639 && 
b[21640] == 21640 && 
b[21641] == 21641 && 
b[21642] == 21642 && 
b[21643] == 21643 && 
b[21644] == 21644 && 
b[21645] == 21645 && 
b[21646] == 21646 && 
b[21647] == 21647 && 
b[21648] == 21648 && 
b[21649] == 21649 && 
b[21650] == 21650 && 
b[21651] == 21651 && 
b[21652] == 21652 && 
b[21653] == 21653 && 
b[21654] == 21654 && 
b[21655] == 21655 && 
b[21656] == 21656 && 
b[21657] == 21657 && 
b[21658] == 21658 && 
b[21659] == 21659 && 
b[21660] == 21660 && 
b[21661] == 21661 && 
b[21662] == 21662 && 
b[21663] == 21663 && 
b[21664] == 21664 && 
b[21665] == 21665 && 
b[21666] == 21666 && 
b[21667] == 21667 && 
b[21668] == 21668 && 
b[21669] == 21669 && 
b[21670] == 21670 && 
b[21671] == 21671 && 
b[21672] == 21672 && 
b[21673] == 21673 && 
b[21674] == 21674 && 
b[21675] == 21675 && 
b[21676] == 21676 && 
b[21677] == 21677 && 
b[21678] == 21678 && 
b[21679] == 21679 && 
b[21680] == 21680 && 
b[21681] == 21681 && 
b[21682] == 21682 && 
b[21683] == 21683 && 
b[21684] == 21684 && 
b[21685] == 21685 && 
b[21686] == 21686 && 
b[21687] == 21687 && 
b[21688] == 21688 && 
b[21689] == 21689 && 
b[21690] == 21690 && 
b[21691] == 21691 && 
b[21692] == 21692 && 
b[21693] == 21693 && 
b[21694] == 21694 && 
b[21695] == 21695 && 
b[21696] == 21696 && 
b[21697] == 21697 && 
b[21698] == 21698 && 
b[21699] == 21699 && 
b[21700] == 21700 && 
b[21701] == 21701 && 
b[21702] == 21702 && 
b[21703] == 21703 && 
b[21704] == 21704 && 
b[21705] == 21705 && 
b[21706] == 21706 && 
b[21707] == 21707 && 
b[21708] == 21708 && 
b[21709] == 21709 && 
b[21710] == 21710 && 
b[21711] == 21711 && 
b[21712] == 21712 && 
b[21713] == 21713 && 
b[21714] == 21714 && 
b[21715] == 21715 && 
b[21716] == 21716 && 
b[21717] == 21717 && 
b[21718] == 21718 && 
b[21719] == 21719 && 
b[21720] == 21720 && 
b[21721] == 21721 && 
b[21722] == 21722 && 
b[21723] == 21723 && 
b[21724] == 21724 && 
b[21725] == 21725 && 
b[21726] == 21726 && 
b[21727] == 21727 && 
b[21728] == 21728 && 
b[21729] == 21729 && 
b[21730] == 21730 && 
b[21731] == 21731 && 
b[21732] == 21732 && 
b[21733] == 21733 && 
b[21734] == 21734 && 
b[21735] == 21735 && 
b[21736] == 21736 && 
b[21737] == 21737 && 
b[21738] == 21738 && 
b[21739] == 21739 && 
b[21740] == 21740 && 
b[21741] == 21741 && 
b[21742] == 21742 && 
b[21743] == 21743 && 
b[21744] == 21744 && 
b[21745] == 21745 && 
b[21746] == 21746 && 
b[21747] == 21747 && 
b[21748] == 21748 && 
b[21749] == 21749 && 
b[21750] == 21750 && 
b[21751] == 21751 && 
b[21752] == 21752 && 
b[21753] == 21753 && 
b[21754] == 21754 && 
b[21755] == 21755 && 
b[21756] == 21756 && 
b[21757] == 21757 && 
b[21758] == 21758 && 
b[21759] == 21759 && 
b[21760] == 21760 && 
b[21761] == 21761 && 
b[21762] == 21762 && 
b[21763] == 21763 && 
b[21764] == 21764 && 
b[21765] == 21765 && 
b[21766] == 21766 && 
b[21767] == 21767 && 
b[21768] == 21768 && 
b[21769] == 21769 && 
b[21770] == 21770 && 
b[21771] == 21771 && 
b[21772] == 21772 && 
b[21773] == 21773 && 
b[21774] == 21774 && 
b[21775] == 21775 && 
b[21776] == 21776 && 
b[21777] == 21777 && 
b[21778] == 21778 && 
b[21779] == 21779 && 
b[21780] == 21780 && 
b[21781] == 21781 && 
b[21782] == 21782 && 
b[21783] == 21783 && 
b[21784] == 21784 && 
b[21785] == 21785 && 
b[21786] == 21786 && 
b[21787] == 21787 && 
b[21788] == 21788 && 
b[21789] == 21789 && 
b[21790] == 21790 && 
b[21791] == 21791 && 
b[21792] == 21792 && 
b[21793] == 21793 && 
b[21794] == 21794 && 
b[21795] == 21795 && 
b[21796] == 21796 && 
b[21797] == 21797 && 
b[21798] == 21798 && 
b[21799] == 21799 && 
b[21800] == 21800 && 
b[21801] == 21801 && 
b[21802] == 21802 && 
b[21803] == 21803 && 
b[21804] == 21804 && 
b[21805] == 21805 && 
b[21806] == 21806 && 
b[21807] == 21807 && 
b[21808] == 21808 && 
b[21809] == 21809 && 
b[21810] == 21810 && 
b[21811] == 21811 && 
b[21812] == 21812 && 
b[21813] == 21813 && 
b[21814] == 21814 && 
b[21815] == 21815 && 
b[21816] == 21816 && 
b[21817] == 21817 && 
b[21818] == 21818 && 
b[21819] == 21819 && 
b[21820] == 21820 && 
b[21821] == 21821 && 
b[21822] == 21822 && 
b[21823] == 21823 && 
b[21824] == 21824 && 
b[21825] == 21825 && 
b[21826] == 21826 && 
b[21827] == 21827 && 
b[21828] == 21828 && 
b[21829] == 21829 && 
b[21830] == 21830 && 
b[21831] == 21831 && 
b[21832] == 21832 && 
b[21833] == 21833 && 
b[21834] == 21834 && 
b[21835] == 21835 && 
b[21836] == 21836 && 
b[21837] == 21837 && 
b[21838] == 21838 && 
b[21839] == 21839 && 
b[21840] == 21840 && 
b[21841] == 21841 && 
b[21842] == 21842 && 
b[21843] == 21843 && 
b[21844] == 21844 && 
b[21845] == 21845 && 
b[21846] == 21846 && 
b[21847] == 21847 && 
b[21848] == 21848 && 
b[21849] == 21849 && 
b[21850] == 21850 && 
b[21851] == 21851 && 
b[21852] == 21852 && 
b[21853] == 21853 && 
b[21854] == 21854 && 
b[21855] == 21855 && 
b[21856] == 21856 && 
b[21857] == 21857 && 
b[21858] == 21858 && 
b[21859] == 21859 && 
b[21860] == 21860 && 
b[21861] == 21861 && 
b[21862] == 21862 && 
b[21863] == 21863 && 
b[21864] == 21864 && 
b[21865] == 21865 && 
b[21866] == 21866 && 
b[21867] == 21867 && 
b[21868] == 21868 && 
b[21869] == 21869 && 
b[21870] == 21870 && 
b[21871] == 21871 && 
b[21872] == 21872 && 
b[21873] == 21873 && 
b[21874] == 21874 && 
b[21875] == 21875 && 
b[21876] == 21876 && 
b[21877] == 21877 && 
b[21878] == 21878 && 
b[21879] == 21879 && 
b[21880] == 21880 && 
b[21881] == 21881 && 
b[21882] == 21882 && 
b[21883] == 21883 && 
b[21884] == 21884 && 
b[21885] == 21885 && 
b[21886] == 21886 && 
b[21887] == 21887 && 
b[21888] == 21888 && 
b[21889] == 21889 && 
b[21890] == 21890 && 
b[21891] == 21891 && 
b[21892] == 21892 && 
b[21893] == 21893 && 
b[21894] == 21894 && 
b[21895] == 21895 && 
b[21896] == 21896 && 
b[21897] == 21897 && 
b[21898] == 21898 && 
b[21899] == 21899 && 
b[21900] == 21900 && 
b[21901] == 21901 && 
b[21902] == 21902 && 
b[21903] == 21903 && 
b[21904] == 21904 && 
b[21905] == 21905 && 
b[21906] == 21906 && 
b[21907] == 21907 && 
b[21908] == 21908 && 
b[21909] == 21909 && 
b[21910] == 21910 && 
b[21911] == 21911 && 
b[21912] == 21912 && 
b[21913] == 21913 && 
b[21914] == 21914 && 
b[21915] == 21915 && 
b[21916] == 21916 && 
b[21917] == 21917 && 
b[21918] == 21918 && 
b[21919] == 21919 && 
b[21920] == 21920 && 
b[21921] == 21921 && 
b[21922] == 21922 && 
b[21923] == 21923 && 
b[21924] == 21924 && 
b[21925] == 21925 && 
b[21926] == 21926 && 
b[21927] == 21927 && 
b[21928] == 21928 && 
b[21929] == 21929 && 
b[21930] == 21930 && 
b[21931] == 21931 && 
b[21932] == 21932 && 
b[21933] == 21933 && 
b[21934] == 21934 && 
b[21935] == 21935 && 
b[21936] == 21936 && 
b[21937] == 21937 && 
b[21938] == 21938 && 
b[21939] == 21939 && 
b[21940] == 21940 && 
b[21941] == 21941 && 
b[21942] == 21942 && 
b[21943] == 21943 && 
b[21944] == 21944 && 
b[21945] == 21945 && 
b[21946] == 21946 && 
b[21947] == 21947 && 
b[21948] == 21948 && 
b[21949] == 21949 && 
b[21950] == 21950 && 
b[21951] == 21951 && 
b[21952] == 21952 && 
b[21953] == 21953 && 
b[21954] == 21954 && 
b[21955] == 21955 && 
b[21956] == 21956 && 
b[21957] == 21957 && 
b[21958] == 21958 && 
b[21959] == 21959 && 
b[21960] == 21960 && 
b[21961] == 21961 && 
b[21962] == 21962 && 
b[21963] == 21963 && 
b[21964] == 21964 && 
b[21965] == 21965 && 
b[21966] == 21966 && 
b[21967] == 21967 && 
b[21968] == 21968 && 
b[21969] == 21969 && 
b[21970] == 21970 && 
b[21971] == 21971 && 
b[21972] == 21972 && 
b[21973] == 21973 && 
b[21974] == 21974 && 
b[21975] == 21975 && 
b[21976] == 21976 && 
b[21977] == 21977 && 
b[21978] == 21978 && 
b[21979] == 21979 && 
b[21980] == 21980 && 
b[21981] == 21981 && 
b[21982] == 21982 && 
b[21983] == 21983 && 
b[21984] == 21984 && 
b[21985] == 21985 && 
b[21986] == 21986 && 
b[21987] == 21987 && 
b[21988] == 21988 && 
b[21989] == 21989 && 
b[21990] == 21990 && 
b[21991] == 21991 && 
b[21992] == 21992 && 
b[21993] == 21993 && 
b[21994] == 21994 && 
b[21995] == 21995 && 
b[21996] == 21996 && 
b[21997] == 21997 && 
b[21998] == 21998 && 
b[21999] == 21999 && 
b[22000] == 22000 && 
b[22001] == 22001 && 
b[22002] == 22002 && 
b[22003] == 22003 && 
b[22004] == 22004 && 
b[22005] == 22005 && 
b[22006] == 22006 && 
b[22007] == 22007 && 
b[22008] == 22008 && 
b[22009] == 22009 && 
b[22010] == 22010 && 
b[22011] == 22011 && 
b[22012] == 22012 && 
b[22013] == 22013 && 
b[22014] == 22014 && 
b[22015] == 22015 && 
b[22016] == 22016 && 
b[22017] == 22017 && 
b[22018] == 22018 && 
b[22019] == 22019 && 
b[22020] == 22020 && 
b[22021] == 22021 && 
b[22022] == 22022 && 
b[22023] == 22023 && 
b[22024] == 22024 && 
b[22025] == 22025 && 
b[22026] == 22026 && 
b[22027] == 22027 && 
b[22028] == 22028 && 
b[22029] == 22029 && 
b[22030] == 22030 && 
b[22031] == 22031 && 
b[22032] == 22032 && 
b[22033] == 22033 && 
b[22034] == 22034 && 
b[22035] == 22035 && 
b[22036] == 22036 && 
b[22037] == 22037 && 
b[22038] == 22038 && 
b[22039] == 22039 && 
b[22040] == 22040 && 
b[22041] == 22041 && 
b[22042] == 22042 && 
b[22043] == 22043 && 
b[22044] == 22044 && 
b[22045] == 22045 && 
b[22046] == 22046 && 
b[22047] == 22047 && 
b[22048] == 22048 && 
b[22049] == 22049 && 
b[22050] == 22050 && 
b[22051] == 22051 && 
b[22052] == 22052 && 
b[22053] == 22053 && 
b[22054] == 22054 && 
b[22055] == 22055 && 
b[22056] == 22056 && 
b[22057] == 22057 && 
b[22058] == 22058 && 
b[22059] == 22059 && 
b[22060] == 22060 && 
b[22061] == 22061 && 
b[22062] == 22062 && 
b[22063] == 22063 && 
b[22064] == 22064 && 
b[22065] == 22065 && 
b[22066] == 22066 && 
b[22067] == 22067 && 
b[22068] == 22068 && 
b[22069] == 22069 && 
b[22070] == 22070 && 
b[22071] == 22071 && 
b[22072] == 22072 && 
b[22073] == 22073 && 
b[22074] == 22074 && 
b[22075] == 22075 && 
b[22076] == 22076 && 
b[22077] == 22077 && 
b[22078] == 22078 && 
b[22079] == 22079 && 
b[22080] == 22080 && 
b[22081] == 22081 && 
b[22082] == 22082 && 
b[22083] == 22083 && 
b[22084] == 22084 && 
b[22085] == 22085 && 
b[22086] == 22086 && 
b[22087] == 22087 && 
b[22088] == 22088 && 
b[22089] == 22089 && 
b[22090] == 22090 && 
b[22091] == 22091 && 
b[22092] == 22092 && 
b[22093] == 22093 && 
b[22094] == 22094 && 
b[22095] == 22095 && 
b[22096] == 22096 && 
b[22097] == 22097 && 
b[22098] == 22098 && 
b[22099] == 22099 && 
b[22100] == 22100 && 
b[22101] == 22101 && 
b[22102] == 22102 && 
b[22103] == 22103 && 
b[22104] == 22104 && 
b[22105] == 22105 && 
b[22106] == 22106 && 
b[22107] == 22107 && 
b[22108] == 22108 && 
b[22109] == 22109 && 
b[22110] == 22110 && 
b[22111] == 22111 && 
b[22112] == 22112 && 
b[22113] == 22113 && 
b[22114] == 22114 && 
b[22115] == 22115 && 
b[22116] == 22116 && 
b[22117] == 22117 && 
b[22118] == 22118 && 
b[22119] == 22119 && 
b[22120] == 22120 && 
b[22121] == 22121 && 
b[22122] == 22122 && 
b[22123] == 22123 && 
b[22124] == 22124 && 
b[22125] == 22125 && 
b[22126] == 22126 && 
b[22127] == 22127 && 
b[22128] == 22128 && 
b[22129] == 22129 && 
b[22130] == 22130 && 
b[22131] == 22131 && 
b[22132] == 22132 && 
b[22133] == 22133 && 
b[22134] == 22134 && 
b[22135] == 22135 && 
b[22136] == 22136 && 
b[22137] == 22137 && 
b[22138] == 22138 && 
b[22139] == 22139 && 
b[22140] == 22140 && 
b[22141] == 22141 && 
b[22142] == 22142 && 
b[22143] == 22143 && 
b[22144] == 22144 && 
b[22145] == 22145 && 
b[22146] == 22146 && 
b[22147] == 22147 && 
b[22148] == 22148 && 
b[22149] == 22149 && 
b[22150] == 22150 && 
b[22151] == 22151 && 
b[22152] == 22152 && 
b[22153] == 22153 && 
b[22154] == 22154 && 
b[22155] == 22155 && 
b[22156] == 22156 && 
b[22157] == 22157 && 
b[22158] == 22158 && 
b[22159] == 22159 && 
b[22160] == 22160 && 
b[22161] == 22161 && 
b[22162] == 22162 && 
b[22163] == 22163 && 
b[22164] == 22164 && 
b[22165] == 22165 && 
b[22166] == 22166 && 
b[22167] == 22167 && 
b[22168] == 22168 && 
b[22169] == 22169 && 
b[22170] == 22170 && 
b[22171] == 22171 && 
b[22172] == 22172 && 
b[22173] == 22173 && 
b[22174] == 22174 && 
b[22175] == 22175 && 
b[22176] == 22176 && 
b[22177] == 22177 && 
b[22178] == 22178 && 
b[22179] == 22179 && 
b[22180] == 22180 && 
b[22181] == 22181 && 
b[22182] == 22182 && 
b[22183] == 22183 && 
b[22184] == 22184 && 
b[22185] == 22185 && 
b[22186] == 22186 && 
b[22187] == 22187 && 
b[22188] == 22188 && 
b[22189] == 22189 && 
b[22190] == 22190 && 
b[22191] == 22191 && 
b[22192] == 22192 && 
b[22193] == 22193 && 
b[22194] == 22194 && 
b[22195] == 22195 && 
b[22196] == 22196 && 
b[22197] == 22197 && 
b[22198] == 22198 && 
b[22199] == 22199 && 
b[22200] == 22200 && 
b[22201] == 22201 && 
b[22202] == 22202 && 
b[22203] == 22203 && 
b[22204] == 22204 && 
b[22205] == 22205 && 
b[22206] == 22206 && 
b[22207] == 22207 && 
b[22208] == 22208 && 
b[22209] == 22209 && 
b[22210] == 22210 && 
b[22211] == 22211 && 
b[22212] == 22212 && 
b[22213] == 22213 && 
b[22214] == 22214 && 
b[22215] == 22215 && 
b[22216] == 22216 && 
b[22217] == 22217 && 
b[22218] == 22218 && 
b[22219] == 22219 && 
b[22220] == 22220 && 
b[22221] == 22221 && 
b[22222] == 22222 && 
b[22223] == 22223 && 
b[22224] == 22224 && 
b[22225] == 22225 && 
b[22226] == 22226 && 
b[22227] == 22227 && 
b[22228] == 22228 && 
b[22229] == 22229 && 
b[22230] == 22230 && 
b[22231] == 22231 && 
b[22232] == 22232 && 
b[22233] == 22233 && 
b[22234] == 22234 && 
b[22235] == 22235 && 
b[22236] == 22236 && 
b[22237] == 22237 && 
b[22238] == 22238 && 
b[22239] == 22239 && 
b[22240] == 22240 && 
b[22241] == 22241 && 
b[22242] == 22242 && 
b[22243] == 22243 && 
b[22244] == 22244 && 
b[22245] == 22245 && 
b[22246] == 22246 && 
b[22247] == 22247 && 
b[22248] == 22248 && 
b[22249] == 22249 && 
b[22250] == 22250 && 
b[22251] == 22251 && 
b[22252] == 22252 && 
b[22253] == 22253 && 
b[22254] == 22254 && 
b[22255] == 22255 && 
b[22256] == 22256 && 
b[22257] == 22257 && 
b[22258] == 22258 && 
b[22259] == 22259 && 
b[22260] == 22260 && 
b[22261] == 22261 && 
b[22262] == 22262 && 
b[22263] == 22263 && 
b[22264] == 22264 && 
b[22265] == 22265 && 
b[22266] == 22266 && 
b[22267] == 22267 && 
b[22268] == 22268 && 
b[22269] == 22269 && 
b[22270] == 22270 && 
b[22271] == 22271 && 
b[22272] == 22272 && 
b[22273] == 22273 && 
b[22274] == 22274 && 
b[22275] == 22275 && 
b[22276] == 22276 && 
b[22277] == 22277 && 
b[22278] == 22278 && 
b[22279] == 22279 && 
b[22280] == 22280 && 
b[22281] == 22281 && 
b[22282] == 22282 && 
b[22283] == 22283 && 
b[22284] == 22284 && 
b[22285] == 22285 && 
b[22286] == 22286 && 
b[22287] == 22287 && 
b[22288] == 22288 && 
b[22289] == 22289 && 
b[22290] == 22290 && 
b[22291] == 22291 && 
b[22292] == 22292 && 
b[22293] == 22293 && 
b[22294] == 22294 && 
b[22295] == 22295 && 
b[22296] == 22296 && 
b[22297] == 22297 && 
b[22298] == 22298 && 
b[22299] == 22299 && 
b[22300] == 22300 && 
b[22301] == 22301 && 
b[22302] == 22302 && 
b[22303] == 22303 && 
b[22304] == 22304 && 
b[22305] == 22305 && 
b[22306] == 22306 && 
b[22307] == 22307 && 
b[22308] == 22308 && 
b[22309] == 22309 && 
b[22310] == 22310 && 
b[22311] == 22311 && 
b[22312] == 22312 && 
b[22313] == 22313 && 
b[22314] == 22314 && 
b[22315] == 22315 && 
b[22316] == 22316 && 
b[22317] == 22317 && 
b[22318] == 22318 && 
b[22319] == 22319 && 
b[22320] == 22320 && 
b[22321] == 22321 && 
b[22322] == 22322 && 
b[22323] == 22323 && 
b[22324] == 22324 && 
b[22325] == 22325 && 
b[22326] == 22326 && 
b[22327] == 22327 && 
b[22328] == 22328 && 
b[22329] == 22329 && 
b[22330] == 22330 && 
b[22331] == 22331 && 
b[22332] == 22332 && 
b[22333] == 22333 && 
b[22334] == 22334 && 
b[22335] == 22335 && 
b[22336] == 22336 && 
b[22337] == 22337 && 
b[22338] == 22338 && 
b[22339] == 22339 && 
b[22340] == 22340 && 
b[22341] == 22341 && 
b[22342] == 22342 && 
b[22343] == 22343 && 
b[22344] == 22344 && 
b[22345] == 22345 && 
b[22346] == 22346 && 
b[22347] == 22347 && 
b[22348] == 22348 && 
b[22349] == 22349 && 
b[22350] == 22350 && 
b[22351] == 22351 && 
b[22352] == 22352 && 
b[22353] == 22353 && 
b[22354] == 22354 && 
b[22355] == 22355 && 
b[22356] == 22356 && 
b[22357] == 22357 && 
b[22358] == 22358 && 
b[22359] == 22359 && 
b[22360] == 22360 && 
b[22361] == 22361 && 
b[22362] == 22362 && 
b[22363] == 22363 && 
b[22364] == 22364 && 
b[22365] == 22365 && 
b[22366] == 22366 && 
b[22367] == 22367 && 
b[22368] == 22368 && 
b[22369] == 22369 && 
b[22370] == 22370 && 
b[22371] == 22371 && 
b[22372] == 22372 && 
b[22373] == 22373 && 
b[22374] == 22374 && 
b[22375] == 22375 && 
b[22376] == 22376 && 
b[22377] == 22377 && 
b[22378] == 22378 && 
b[22379] == 22379 && 
b[22380] == 22380 && 
b[22381] == 22381 && 
b[22382] == 22382 && 
b[22383] == 22383 && 
b[22384] == 22384 && 
b[22385] == 22385 && 
b[22386] == 22386 && 
b[22387] == 22387 && 
b[22388] == 22388 && 
b[22389] == 22389 && 
b[22390] == 22390 && 
b[22391] == 22391 && 
b[22392] == 22392 && 
b[22393] == 22393 && 
b[22394] == 22394 && 
b[22395] == 22395 && 
b[22396] == 22396 && 
b[22397] == 22397 && 
b[22398] == 22398 && 
b[22399] == 22399 && 
b[22400] == 22400 && 
b[22401] == 22401 && 
b[22402] == 22402 && 
b[22403] == 22403 && 
b[22404] == 22404 && 
b[22405] == 22405 && 
b[22406] == 22406 && 
b[22407] == 22407 && 
b[22408] == 22408 && 
b[22409] == 22409 && 
b[22410] == 22410 && 
b[22411] == 22411 && 
b[22412] == 22412 && 
b[22413] == 22413 && 
b[22414] == 22414 && 
b[22415] == 22415 && 
b[22416] == 22416 && 
b[22417] == 22417 && 
b[22418] == 22418 && 
b[22419] == 22419 && 
b[22420] == 22420 && 
b[22421] == 22421 && 
b[22422] == 22422 && 
b[22423] == 22423 && 
b[22424] == 22424 && 
b[22425] == 22425 && 
b[22426] == 22426 && 
b[22427] == 22427 && 
b[22428] == 22428 && 
b[22429] == 22429 && 
b[22430] == 22430 && 
b[22431] == 22431 && 
b[22432] == 22432 && 
b[22433] == 22433 && 
b[22434] == 22434 && 
b[22435] == 22435 && 
b[22436] == 22436 && 
b[22437] == 22437 && 
b[22438] == 22438 && 
b[22439] == 22439 && 
b[22440] == 22440 && 
b[22441] == 22441 && 
b[22442] == 22442 && 
b[22443] == 22443 && 
b[22444] == 22444 && 
b[22445] == 22445 && 
b[22446] == 22446 && 
b[22447] == 22447 && 
b[22448] == 22448 && 
b[22449] == 22449 && 
b[22450] == 22450 && 
b[22451] == 22451 && 
b[22452] == 22452 && 
b[22453] == 22453 && 
b[22454] == 22454 && 
b[22455] == 22455 && 
b[22456] == 22456 && 
b[22457] == 22457 && 
b[22458] == 22458 && 
b[22459] == 22459 && 
b[22460] == 22460 && 
b[22461] == 22461 && 
b[22462] == 22462 && 
b[22463] == 22463 && 
b[22464] == 22464 && 
b[22465] == 22465 && 
b[22466] == 22466 && 
b[22467] == 22467 && 
b[22468] == 22468 && 
b[22469] == 22469 && 
b[22470] == 22470 && 
b[22471] == 22471 && 
b[22472] == 22472 && 
b[22473] == 22473 && 
b[22474] == 22474 && 
b[22475] == 22475 && 
b[22476] == 22476 && 
b[22477] == 22477 && 
b[22478] == 22478 && 
b[22479] == 22479 && 
b[22480] == 22480 && 
b[22481] == 22481 && 
b[22482] == 22482 && 
b[22483] == 22483 && 
b[22484] == 22484 && 
b[22485] == 22485 && 
b[22486] == 22486 && 
b[22487] == 22487 && 
b[22488] == 22488 && 
b[22489] == 22489 && 
b[22490] == 22490 && 
b[22491] == 22491 && 
b[22492] == 22492 && 
b[22493] == 22493 && 
b[22494] == 22494 && 
b[22495] == 22495 && 
b[22496] == 22496 && 
b[22497] == 22497 && 
b[22498] == 22498 && 
b[22499] == 22499 && 
b[22500] == 22500 && 
b[22501] == 22501 && 
b[22502] == 22502 && 
b[22503] == 22503 && 
b[22504] == 22504 && 
b[22505] == 22505 && 
b[22506] == 22506 && 
b[22507] == 22507 && 
b[22508] == 22508 && 
b[22509] == 22509 && 
b[22510] == 22510 && 
b[22511] == 22511 && 
b[22512] == 22512 && 
b[22513] == 22513 && 
b[22514] == 22514 && 
b[22515] == 22515 && 
b[22516] == 22516 && 
b[22517] == 22517 && 
b[22518] == 22518 && 
b[22519] == 22519 && 
b[22520] == 22520 && 
b[22521] == 22521 && 
b[22522] == 22522 && 
b[22523] == 22523 && 
b[22524] == 22524 && 
b[22525] == 22525 && 
b[22526] == 22526 && 
b[22527] == 22527 && 
b[22528] == 22528 && 
b[22529] == 22529 && 
b[22530] == 22530 && 
b[22531] == 22531 && 
b[22532] == 22532 && 
b[22533] == 22533 && 
b[22534] == 22534 && 
b[22535] == 22535 && 
b[22536] == 22536 && 
b[22537] == 22537 && 
b[22538] == 22538 && 
b[22539] == 22539 && 
b[22540] == 22540 && 
b[22541] == 22541 && 
b[22542] == 22542 && 
b[22543] == 22543 && 
b[22544] == 22544 && 
b[22545] == 22545 && 
b[22546] == 22546 && 
b[22547] == 22547 && 
b[22548] == 22548 && 
b[22549] == 22549 && 
b[22550] == 22550 && 
b[22551] == 22551 && 
b[22552] == 22552 && 
b[22553] == 22553 && 
b[22554] == 22554 && 
b[22555] == 22555 && 
b[22556] == 22556 && 
b[22557] == 22557 && 
b[22558] == 22558 && 
b[22559] == 22559 && 
b[22560] == 22560 && 
b[22561] == 22561 && 
b[22562] == 22562 && 
b[22563] == 22563 && 
b[22564] == 22564 && 
b[22565] == 22565 && 
b[22566] == 22566 && 
b[22567] == 22567 && 
b[22568] == 22568 && 
b[22569] == 22569 && 
b[22570] == 22570 && 
b[22571] == 22571 && 
b[22572] == 22572 && 
b[22573] == 22573 && 
b[22574] == 22574 && 
b[22575] == 22575 && 
b[22576] == 22576 && 
b[22577] == 22577 && 
b[22578] == 22578 && 
b[22579] == 22579 && 
b[22580] == 22580 && 
b[22581] == 22581 && 
b[22582] == 22582 && 
b[22583] == 22583 && 
b[22584] == 22584 && 
b[22585] == 22585 && 
b[22586] == 22586 && 
b[22587] == 22587 && 
b[22588] == 22588 && 
b[22589] == 22589 && 
b[22590] == 22590 && 
b[22591] == 22591 && 
b[22592] == 22592 && 
b[22593] == 22593 && 
b[22594] == 22594 && 
b[22595] == 22595 && 
b[22596] == 22596 && 
b[22597] == 22597 && 
b[22598] == 22598 && 
b[22599] == 22599 && 
b[22600] == 22600 && 
b[22601] == 22601 && 
b[22602] == 22602 && 
b[22603] == 22603 && 
b[22604] == 22604 && 
b[22605] == 22605 && 
b[22606] == 22606 && 
b[22607] == 22607 && 
b[22608] == 22608 && 
b[22609] == 22609 && 
b[22610] == 22610 && 
b[22611] == 22611 && 
b[22612] == 22612 && 
b[22613] == 22613 && 
b[22614] == 22614 && 
b[22615] == 22615 && 
b[22616] == 22616 && 
b[22617] == 22617 && 
b[22618] == 22618 && 
b[22619] == 22619 && 
b[22620] == 22620 && 
b[22621] == 22621 && 
b[22622] == 22622 && 
b[22623] == 22623 && 
b[22624] == 22624 && 
b[22625] == 22625 && 
b[22626] == 22626 && 
b[22627] == 22627 && 
b[22628] == 22628 && 
b[22629] == 22629 && 
b[22630] == 22630 && 
b[22631] == 22631 && 
b[22632] == 22632 && 
b[22633] == 22633 && 
b[22634] == 22634 && 
b[22635] == 22635 && 
b[22636] == 22636 && 
b[22637] == 22637 && 
b[22638] == 22638 && 
b[22639] == 22639 && 
b[22640] == 22640 && 
b[22641] == 22641 && 
b[22642] == 22642 && 
b[22643] == 22643 && 
b[22644] == 22644 && 
b[22645] == 22645 && 
b[22646] == 22646 && 
b[22647] == 22647 && 
b[22648] == 22648 && 
b[22649] == 22649 && 
b[22650] == 22650 && 
b[22651] == 22651 && 
b[22652] == 22652 && 
b[22653] == 22653 && 
b[22654] == 22654 && 
b[22655] == 22655 && 
b[22656] == 22656 && 
b[22657] == 22657 && 
b[22658] == 22658 && 
b[22659] == 22659 && 
b[22660] == 22660 && 
b[22661] == 22661 && 
b[22662] == 22662 && 
b[22663] == 22663 && 
b[22664] == 22664 && 
b[22665] == 22665 && 
b[22666] == 22666 && 
b[22667] == 22667 && 
b[22668] == 22668 && 
b[22669] == 22669 && 
b[22670] == 22670 && 
b[22671] == 22671 && 
b[22672] == 22672 && 
b[22673] == 22673 && 
b[22674] == 22674 && 
b[22675] == 22675 && 
b[22676] == 22676 && 
b[22677] == 22677 && 
b[22678] == 22678 && 
b[22679] == 22679 && 
b[22680] == 22680 && 
b[22681] == 22681 && 
b[22682] == 22682 && 
b[22683] == 22683 && 
b[22684] == 22684 && 
b[22685] == 22685 && 
b[22686] == 22686 && 
b[22687] == 22687 && 
b[22688] == 22688 && 
b[22689] == 22689 && 
b[22690] == 22690 && 
b[22691] == 22691 && 
b[22692] == 22692 && 
b[22693] == 22693 && 
b[22694] == 22694 && 
b[22695] == 22695 && 
b[22696] == 22696 && 
b[22697] == 22697 && 
b[22698] == 22698 && 
b[22699] == 22699 && 
b[22700] == 22700 && 
b[22701] == 22701 && 
b[22702] == 22702 && 
b[22703] == 22703 && 
b[22704] == 22704 && 
b[22705] == 22705 && 
b[22706] == 22706 && 
b[22707] == 22707 && 
b[22708] == 22708 && 
b[22709] == 22709 && 
b[22710] == 22710 && 
b[22711] == 22711 && 
b[22712] == 22712 && 
b[22713] == 22713 && 
b[22714] == 22714 && 
b[22715] == 22715 && 
b[22716] == 22716 && 
b[22717] == 22717 && 
b[22718] == 22718 && 
b[22719] == 22719 && 
b[22720] == 22720 && 
b[22721] == 22721 && 
b[22722] == 22722 && 
b[22723] == 22723 && 
b[22724] == 22724 && 
b[22725] == 22725 && 
b[22726] == 22726 && 
b[22727] == 22727 && 
b[22728] == 22728 && 
b[22729] == 22729 && 
b[22730] == 22730 && 
b[22731] == 22731 && 
b[22732] == 22732 && 
b[22733] == 22733 && 
b[22734] == 22734 && 
b[22735] == 22735 && 
b[22736] == 22736 && 
b[22737] == 22737 && 
b[22738] == 22738 && 
b[22739] == 22739 && 
b[22740] == 22740 && 
b[22741] == 22741 && 
b[22742] == 22742 && 
b[22743] == 22743 && 
b[22744] == 22744 && 
b[22745] == 22745 && 
b[22746] == 22746 && 
b[22747] == 22747 && 
b[22748] == 22748 && 
b[22749] == 22749 && 
b[22750] == 22750 && 
b[22751] == 22751 && 
b[22752] == 22752 && 
b[22753] == 22753 && 
b[22754] == 22754 && 
b[22755] == 22755 && 
b[22756] == 22756 && 
b[22757] == 22757 && 
b[22758] == 22758 && 
b[22759] == 22759 && 
b[22760] == 22760 && 
b[22761] == 22761 && 
b[22762] == 22762 && 
b[22763] == 22763 && 
b[22764] == 22764 && 
b[22765] == 22765 && 
b[22766] == 22766 && 
b[22767] == 22767 && 
b[22768] == 22768 && 
b[22769] == 22769 && 
b[22770] == 22770 && 
b[22771] == 22771 && 
b[22772] == 22772 && 
b[22773] == 22773 && 
b[22774] == 22774 && 
b[22775] == 22775 && 
b[22776] == 22776 && 
b[22777] == 22777 && 
b[22778] == 22778 && 
b[22779] == 22779 && 
b[22780] == 22780 && 
b[22781] == 22781 && 
b[22782] == 22782 && 
b[22783] == 22783 && 
b[22784] == 22784 && 
b[22785] == 22785 && 
b[22786] == 22786 && 
b[22787] == 22787 && 
b[22788] == 22788 && 
b[22789] == 22789 && 
b[22790] == 22790 && 
b[22791] == 22791 && 
b[22792] == 22792 && 
b[22793] == 22793 && 
b[22794] == 22794 && 
b[22795] == 22795 && 
b[22796] == 22796 && 
b[22797] == 22797 && 
b[22798] == 22798 && 
b[22799] == 22799 && 
b[22800] == 22800 && 
b[22801] == 22801 && 
b[22802] == 22802 && 
b[22803] == 22803 && 
b[22804] == 22804 && 
b[22805] == 22805 && 
b[22806] == 22806 && 
b[22807] == 22807 && 
b[22808] == 22808 && 
b[22809] == 22809 && 
b[22810] == 22810 && 
b[22811] == 22811 && 
b[22812] == 22812 && 
b[22813] == 22813 && 
b[22814] == 22814 && 
b[22815] == 22815 && 
b[22816] == 22816 && 
b[22817] == 22817 && 
b[22818] == 22818 && 
b[22819] == 22819 && 
b[22820] == 22820 && 
b[22821] == 22821 && 
b[22822] == 22822 && 
b[22823] == 22823 && 
b[22824] == 22824 && 
b[22825] == 22825 && 
b[22826] == 22826 && 
b[22827] == 22827 && 
b[22828] == 22828 && 
b[22829] == 22829 && 
b[22830] == 22830 && 
b[22831] == 22831 && 
b[22832] == 22832 && 
b[22833] == 22833 && 
b[22834] == 22834 && 
b[22835] == 22835 && 
b[22836] == 22836 && 
b[22837] == 22837 && 
b[22838] == 22838 && 
b[22839] == 22839 && 
b[22840] == 22840 && 
b[22841] == 22841 && 
b[22842] == 22842 && 
b[22843] == 22843 && 
b[22844] == 22844 && 
b[22845] == 22845 && 
b[22846] == 22846 && 
b[22847] == 22847 && 
b[22848] == 22848 && 
b[22849] == 22849 && 
b[22850] == 22850 && 
b[22851] == 22851 && 
b[22852] == 22852 && 
b[22853] == 22853 && 
b[22854] == 22854 && 
b[22855] == 22855 && 
b[22856] == 22856 && 
b[22857] == 22857 && 
b[22858] == 22858 && 
b[22859] == 22859 && 
b[22860] == 22860 && 
b[22861] == 22861 && 
b[22862] == 22862 && 
b[22863] == 22863 && 
b[22864] == 22864 && 
b[22865] == 22865 && 
b[22866] == 22866 && 
b[22867] == 22867 && 
b[22868] == 22868 && 
b[22869] == 22869 && 
b[22870] == 22870 && 
b[22871] == 22871 && 
b[22872] == 22872 && 
b[22873] == 22873 && 
b[22874] == 22874 && 
b[22875] == 22875 && 
b[22876] == 22876 && 
b[22877] == 22877 && 
b[22878] == 22878 && 
b[22879] == 22879 && 
b[22880] == 22880 && 
b[22881] == 22881 && 
b[22882] == 22882 && 
b[22883] == 22883 && 
b[22884] == 22884 && 
b[22885] == 22885 && 
b[22886] == 22886 && 
b[22887] == 22887 && 
b[22888] == 22888 && 
b[22889] == 22889 && 
b[22890] == 22890 && 
b[22891] == 22891 && 
b[22892] == 22892 && 
b[22893] == 22893 && 
b[22894] == 22894 && 
b[22895] == 22895 && 
b[22896] == 22896 && 
b[22897] == 22897 && 
b[22898] == 22898 && 
b[22899] == 22899 && 
b[22900] == 22900 && 
b[22901] == 22901 && 
b[22902] == 22902 && 
b[22903] == 22903 && 
b[22904] == 22904 && 
b[22905] == 22905 && 
b[22906] == 22906 && 
b[22907] == 22907 && 
b[22908] == 22908 && 
b[22909] == 22909 && 
b[22910] == 22910 && 
b[22911] == 22911 && 
b[22912] == 22912 && 
b[22913] == 22913 && 
b[22914] == 22914 && 
b[22915] == 22915 && 
b[22916] == 22916 && 
b[22917] == 22917 && 
b[22918] == 22918 && 
b[22919] == 22919 && 
b[22920] == 22920 && 
b[22921] == 22921 && 
b[22922] == 22922 && 
b[22923] == 22923 && 
b[22924] == 22924 && 
b[22925] == 22925 && 
b[22926] == 22926 && 
b[22927] == 22927 && 
b[22928] == 22928 && 
b[22929] == 22929 && 
b[22930] == 22930 && 
b[22931] == 22931 && 
b[22932] == 22932 && 
b[22933] == 22933 && 
b[22934] == 22934 && 
b[22935] == 22935 && 
b[22936] == 22936 && 
b[22937] == 22937 && 
b[22938] == 22938 && 
b[22939] == 22939 && 
b[22940] == 22940 && 
b[22941] == 22941 && 
b[22942] == 22942 && 
b[22943] == 22943 && 
b[22944] == 22944 && 
b[22945] == 22945 && 
b[22946] == 22946 && 
b[22947] == 22947 && 
b[22948] == 22948 && 
b[22949] == 22949 && 
b[22950] == 22950 && 
b[22951] == 22951 && 
b[22952] == 22952 && 
b[22953] == 22953 && 
b[22954] == 22954 && 
b[22955] == 22955 && 
b[22956] == 22956 && 
b[22957] == 22957 && 
b[22958] == 22958 && 
b[22959] == 22959 && 
b[22960] == 22960 && 
b[22961] == 22961 && 
b[22962] == 22962 && 
b[22963] == 22963 && 
b[22964] == 22964 && 
b[22965] == 22965 && 
b[22966] == 22966 && 
b[22967] == 22967 && 
b[22968] == 22968 && 
b[22969] == 22969 && 
b[22970] == 22970 && 
b[22971] == 22971 && 
b[22972] == 22972 && 
b[22973] == 22973 && 
b[22974] == 22974 && 
b[22975] == 22975 && 
b[22976] == 22976 && 
b[22977] == 22977 && 
b[22978] == 22978 && 
b[22979] == 22979 && 
b[22980] == 22980 && 
b[22981] == 22981 && 
b[22982] == 22982 && 
b[22983] == 22983 && 
b[22984] == 22984 && 
b[22985] == 22985 && 
b[22986] == 22986 && 
b[22987] == 22987 && 
b[22988] == 22988 && 
b[22989] == 22989 && 
b[22990] == 22990 && 
b[22991] == 22991 && 
b[22992] == 22992 && 
b[22993] == 22993 && 
b[22994] == 22994 && 
b[22995] == 22995 && 
b[22996] == 22996 && 
b[22997] == 22997 && 
b[22998] == 22998 && 
b[22999] == 22999 && 
b[23000] == 23000 && 
b[23001] == 23001 && 
b[23002] == 23002 && 
b[23003] == 23003 && 
b[23004] == 23004 && 
b[23005] == 23005 && 
b[23006] == 23006 && 
b[23007] == 23007 && 
b[23008] == 23008 && 
b[23009] == 23009 && 
b[23010] == 23010 && 
b[23011] == 23011 && 
b[23012] == 23012 && 
b[23013] == 23013 && 
b[23014] == 23014 && 
b[23015] == 23015 && 
b[23016] == 23016 && 
b[23017] == 23017 && 
b[23018] == 23018 && 
b[23019] == 23019 && 
b[23020] == 23020 && 
b[23021] == 23021 && 
b[23022] == 23022 && 
b[23023] == 23023 && 
b[23024] == 23024 && 
b[23025] == 23025 && 
b[23026] == 23026 && 
b[23027] == 23027 && 
b[23028] == 23028 && 
b[23029] == 23029 && 
b[23030] == 23030 && 
b[23031] == 23031 && 
b[23032] == 23032 && 
b[23033] == 23033 && 
b[23034] == 23034 && 
b[23035] == 23035 && 
b[23036] == 23036 && 
b[23037] == 23037 && 
b[23038] == 23038 && 
b[23039] == 23039 && 
b[23040] == 23040 && 
b[23041] == 23041 && 
b[23042] == 23042 && 
b[23043] == 23043 && 
b[23044] == 23044 && 
b[23045] == 23045 && 
b[23046] == 23046 && 
b[23047] == 23047 && 
b[23048] == 23048 && 
b[23049] == 23049 && 
b[23050] == 23050 && 
b[23051] == 23051 && 
b[23052] == 23052 && 
b[23053] == 23053 && 
b[23054] == 23054 && 
b[23055] == 23055 && 
b[23056] == 23056 && 
b[23057] == 23057 && 
b[23058] == 23058 && 
b[23059] == 23059 && 
b[23060] == 23060 && 
b[23061] == 23061 && 
b[23062] == 23062 && 
b[23063] == 23063 && 
b[23064] == 23064 && 
b[23065] == 23065 && 
b[23066] == 23066 && 
b[23067] == 23067 && 
b[23068] == 23068 && 
b[23069] == 23069 && 
b[23070] == 23070 && 
b[23071] == 23071 && 
b[23072] == 23072 && 
b[23073] == 23073 && 
b[23074] == 23074 && 
b[23075] == 23075 && 
b[23076] == 23076 && 
b[23077] == 23077 && 
b[23078] == 23078 && 
b[23079] == 23079 && 
b[23080] == 23080 && 
b[23081] == 23081 && 
b[23082] == 23082 && 
b[23083] == 23083 && 
b[23084] == 23084 && 
b[23085] == 23085 && 
b[23086] == 23086 && 
b[23087] == 23087 && 
b[23088] == 23088 && 
b[23089] == 23089 && 
b[23090] == 23090 && 
b[23091] == 23091 && 
b[23092] == 23092 && 
b[23093] == 23093 && 
b[23094] == 23094 && 
b[23095] == 23095 && 
b[23096] == 23096 && 
b[23097] == 23097 && 
b[23098] == 23098 && 
b[23099] == 23099 && 
b[23100] == 23100 && 
b[23101] == 23101 && 
b[23102] == 23102 && 
b[23103] == 23103 && 
b[23104] == 23104 && 
b[23105] == 23105 && 
b[23106] == 23106 && 
b[23107] == 23107 && 
b[23108] == 23108 && 
b[23109] == 23109 && 
b[23110] == 23110 && 
b[23111] == 23111 && 
b[23112] == 23112 && 
b[23113] == 23113 && 
b[23114] == 23114 && 
b[23115] == 23115 && 
b[23116] == 23116 && 
b[23117] == 23117 && 
b[23118] == 23118 && 
b[23119] == 23119 && 
b[23120] == 23120 && 
b[23121] == 23121 && 
b[23122] == 23122 && 
b[23123] == 23123 && 
b[23124] == 23124 && 
b[23125] == 23125 && 
b[23126] == 23126 && 
b[23127] == 23127 && 
b[23128] == 23128 && 
b[23129] == 23129 && 
b[23130] == 23130 && 
b[23131] == 23131 && 
b[23132] == 23132 && 
b[23133] == 23133 && 
b[23134] == 23134 && 
b[23135] == 23135 && 
b[23136] == 23136 && 
b[23137] == 23137 && 
b[23138] == 23138 && 
b[23139] == 23139 && 
b[23140] == 23140 && 
b[23141] == 23141 && 
b[23142] == 23142 && 
b[23143] == 23143 && 
b[23144] == 23144 && 
b[23145] == 23145 && 
b[23146] == 23146 && 
b[23147] == 23147 && 
b[23148] == 23148 && 
b[23149] == 23149 && 
b[23150] == 23150 && 
b[23151] == 23151 && 
b[23152] == 23152 && 
b[23153] == 23153 && 
b[23154] == 23154 && 
b[23155] == 23155 && 
b[23156] == 23156 && 
b[23157] == 23157 && 
b[23158] == 23158 && 
b[23159] == 23159 && 
b[23160] == 23160 && 
b[23161] == 23161 && 
b[23162] == 23162 && 
b[23163] == 23163 && 
b[23164] == 23164 && 
b[23165] == 23165 && 
b[23166] == 23166 && 
b[23167] == 23167 && 
b[23168] == 23168 && 
b[23169] == 23169 && 
b[23170] == 23170 && 
b[23171] == 23171 && 
b[23172] == 23172 && 
b[23173] == 23173 && 
b[23174] == 23174 && 
b[23175] == 23175 && 
b[23176] == 23176 && 
b[23177] == 23177 && 
b[23178] == 23178 && 
b[23179] == 23179 && 
b[23180] == 23180 && 
b[23181] == 23181 && 
b[23182] == 23182 && 
b[23183] == 23183 && 
b[23184] == 23184 && 
b[23185] == 23185 && 
b[23186] == 23186 && 
b[23187] == 23187 && 
b[23188] == 23188 && 
b[23189] == 23189 && 
b[23190] == 23190 && 
b[23191] == 23191 && 
b[23192] == 23192 && 
b[23193] == 23193 && 
b[23194] == 23194 && 
b[23195] == 23195 && 
b[23196] == 23196 && 
b[23197] == 23197 && 
b[23198] == 23198 && 
b[23199] == 23199 && 
b[23200] == 23200 && 
b[23201] == 23201 && 
b[23202] == 23202 && 
b[23203] == 23203 && 
b[23204] == 23204 && 
b[23205] == 23205 && 
b[23206] == 23206 && 
b[23207] == 23207 && 
b[23208] == 23208 && 
b[23209] == 23209 && 
b[23210] == 23210 && 
b[23211] == 23211 && 
b[23212] == 23212 && 
b[23213] == 23213 && 
b[23214] == 23214 && 
b[23215] == 23215 && 
b[23216] == 23216 && 
b[23217] == 23217 && 
b[23218] == 23218 && 
b[23219] == 23219 && 
b[23220] == 23220 && 
b[23221] == 23221 && 
b[23222] == 23222 && 
b[23223] == 23223 && 
b[23224] == 23224 && 
b[23225] == 23225 && 
b[23226] == 23226 && 
b[23227] == 23227 && 
b[23228] == 23228 && 
b[23229] == 23229 && 
b[23230] == 23230 && 
b[23231] == 23231 && 
b[23232] == 23232 && 
b[23233] == 23233 && 
b[23234] == 23234 && 
b[23235] == 23235 && 
b[23236] == 23236 && 
b[23237] == 23237 && 
b[23238] == 23238 && 
b[23239] == 23239 && 
b[23240] == 23240 && 
b[23241] == 23241 && 
b[23242] == 23242 && 
b[23243] == 23243 && 
b[23244] == 23244 && 
b[23245] == 23245 && 
b[23246] == 23246 && 
b[23247] == 23247 && 
b[23248] == 23248 && 
b[23249] == 23249 && 
b[23250] == 23250 && 
b[23251] == 23251 && 
b[23252] == 23252 && 
b[23253] == 23253 && 
b[23254] == 23254 && 
b[23255] == 23255 && 
b[23256] == 23256 && 
b[23257] == 23257 && 
b[23258] == 23258 && 
b[23259] == 23259 && 
b[23260] == 23260 && 
b[23261] == 23261 && 
b[23262] == 23262 && 
b[23263] == 23263 && 
b[23264] == 23264 && 
b[23265] == 23265 && 
b[23266] == 23266 && 
b[23267] == 23267 && 
b[23268] == 23268 && 
b[23269] == 23269 && 
b[23270] == 23270 && 
b[23271] == 23271 && 
b[23272] == 23272 && 
b[23273] == 23273 && 
b[23274] == 23274 && 
b[23275] == 23275 && 
b[23276] == 23276 && 
b[23277] == 23277 && 
b[23278] == 23278 && 
b[23279] == 23279 && 
b[23280] == 23280 && 
b[23281] == 23281 && 
b[23282] == 23282 && 
b[23283] == 23283 && 
b[23284] == 23284 && 
b[23285] == 23285 && 
b[23286] == 23286 && 
b[23287] == 23287 && 
b[23288] == 23288 && 
b[23289] == 23289 && 
b[23290] == 23290 && 
b[23291] == 23291 && 
b[23292] == 23292 && 
b[23293] == 23293 && 
b[23294] == 23294 && 
b[23295] == 23295 && 
b[23296] == 23296 && 
b[23297] == 23297 && 
b[23298] == 23298 && 
b[23299] == 23299 && 
b[23300] == 23300 && 
b[23301] == 23301 && 
b[23302] == 23302 && 
b[23303] == 23303 && 
b[23304] == 23304 && 
b[23305] == 23305 && 
b[23306] == 23306 && 
b[23307] == 23307 && 
b[23308] == 23308 && 
b[23309] == 23309 && 
b[23310] == 23310 && 
b[23311] == 23311 && 
b[23312] == 23312 && 
b[23313] == 23313 && 
b[23314] == 23314 && 
b[23315] == 23315 && 
b[23316] == 23316 && 
b[23317] == 23317 && 
b[23318] == 23318 && 
b[23319] == 23319 && 
b[23320] == 23320 && 
b[23321] == 23321 && 
b[23322] == 23322 && 
b[23323] == 23323 && 
b[23324] == 23324 && 
b[23325] == 23325 && 
b[23326] == 23326 && 
b[23327] == 23327 && 
b[23328] == 23328 && 
b[23329] == 23329 && 
b[23330] == 23330 && 
b[23331] == 23331 && 
b[23332] == 23332 && 
b[23333] == 23333 && 
b[23334] == 23334 && 
b[23335] == 23335 && 
b[23336] == 23336 && 
b[23337] == 23337 && 
b[23338] == 23338 && 
b[23339] == 23339 && 
b[23340] == 23340 && 
b[23341] == 23341 && 
b[23342] == 23342 && 
b[23343] == 23343 && 
b[23344] == 23344 && 
b[23345] == 23345 && 
b[23346] == 23346 && 
b[23347] == 23347 && 
b[23348] == 23348 && 
b[23349] == 23349 && 
b[23350] == 23350 && 
b[23351] == 23351 && 
b[23352] == 23352 && 
b[23353] == 23353 && 
b[23354] == 23354 && 
b[23355] == 23355 && 
b[23356] == 23356 && 
b[23357] == 23357 && 
b[23358] == 23358 && 
b[23359] == 23359 && 
b[23360] == 23360 && 
b[23361] == 23361 && 
b[23362] == 23362 && 
b[23363] == 23363 && 
b[23364] == 23364 && 
b[23365] == 23365 && 
b[23366] == 23366 && 
b[23367] == 23367 && 
b[23368] == 23368 && 
b[23369] == 23369 && 
b[23370] == 23370 && 
b[23371] == 23371 && 
b[23372] == 23372 && 
b[23373] == 23373 && 
b[23374] == 23374 && 
b[23375] == 23375 && 
b[23376] == 23376 && 
b[23377] == 23377 && 
b[23378] == 23378 && 
b[23379] == 23379 && 
b[23380] == 23380 && 
b[23381] == 23381 && 
b[23382] == 23382 && 
b[23383] == 23383 && 
b[23384] == 23384 && 
b[23385] == 23385 && 
b[23386] == 23386 && 
b[23387] == 23387 && 
b[23388] == 23388 && 
b[23389] == 23389 && 
b[23390] == 23390 && 
b[23391] == 23391 && 
b[23392] == 23392 && 
b[23393] == 23393 && 
b[23394] == 23394 && 
b[23395] == 23395 && 
b[23396] == 23396 && 
b[23397] == 23397 && 
b[23398] == 23398 && 
b[23399] == 23399 && 
b[23400] == 23400 && 
b[23401] == 23401 && 
b[23402] == 23402 && 
b[23403] == 23403 && 
b[23404] == 23404 && 
b[23405] == 23405 && 
b[23406] == 23406 && 
b[23407] == 23407 && 
b[23408] == 23408 && 
b[23409] == 23409 && 
b[23410] == 23410 && 
b[23411] == 23411 && 
b[23412] == 23412 && 
b[23413] == 23413 && 
b[23414] == 23414 && 
b[23415] == 23415 && 
b[23416] == 23416 && 
b[23417] == 23417 && 
b[23418] == 23418 && 
b[23419] == 23419 && 
b[23420] == 23420 && 
b[23421] == 23421 && 
b[23422] == 23422 && 
b[23423] == 23423 && 
b[23424] == 23424 && 
b[23425] == 23425 && 
b[23426] == 23426 && 
b[23427] == 23427 && 
b[23428] == 23428 && 
b[23429] == 23429 && 
b[23430] == 23430 && 
b[23431] == 23431 && 
b[23432] == 23432 && 
b[23433] == 23433 && 
b[23434] == 23434 && 
b[23435] == 23435 && 
b[23436] == 23436 && 
b[23437] == 23437 && 
b[23438] == 23438 && 
b[23439] == 23439 && 
b[23440] == 23440 && 
b[23441] == 23441 && 
b[23442] == 23442 && 
b[23443] == 23443 && 
b[23444] == 23444 && 
b[23445] == 23445 && 
b[23446] == 23446 && 
b[23447] == 23447 && 
b[23448] == 23448 && 
b[23449] == 23449 && 
b[23450] == 23450 && 
b[23451] == 23451 && 
b[23452] == 23452 && 
b[23453] == 23453 && 
b[23454] == 23454 && 
b[23455] == 23455 && 
b[23456] == 23456 && 
b[23457] == 23457 && 
b[23458] == 23458 && 
b[23459] == 23459 && 
b[23460] == 23460 && 
b[23461] == 23461 && 
b[23462] == 23462 && 
b[23463] == 23463 && 
b[23464] == 23464 && 
b[23465] == 23465 && 
b[23466] == 23466 && 
b[23467] == 23467 && 
b[23468] == 23468 && 
b[23469] == 23469 && 
b[23470] == 23470 && 
b[23471] == 23471 && 
b[23472] == 23472 && 
b[23473] == 23473 && 
b[23474] == 23474 && 
b[23475] == 23475 && 
b[23476] == 23476 && 
b[23477] == 23477 && 
b[23478] == 23478 && 
b[23479] == 23479 && 
b[23480] == 23480 && 
b[23481] == 23481 && 
b[23482] == 23482 && 
b[23483] == 23483 && 
b[23484] == 23484 && 
b[23485] == 23485 && 
b[23486] == 23486 && 
b[23487] == 23487 && 
b[23488] == 23488 && 
b[23489] == 23489 && 
b[23490] == 23490 && 
b[23491] == 23491 && 
b[23492] == 23492 && 
b[23493] == 23493 && 
b[23494] == 23494 && 
b[23495] == 23495 && 
b[23496] == 23496 && 
b[23497] == 23497 && 
b[23498] == 23498 && 
b[23499] == 23499 && 
b[23500] == 23500 && 
b[23501] == 23501 && 
b[23502] == 23502 && 
b[23503] == 23503 && 
b[23504] == 23504 && 
b[23505] == 23505 && 
b[23506] == 23506 && 
b[23507] == 23507 && 
b[23508] == 23508 && 
b[23509] == 23509 && 
b[23510] == 23510 && 
b[23511] == 23511 && 
b[23512] == 23512 && 
b[23513] == 23513 && 
b[23514] == 23514 && 
b[23515] == 23515 && 
b[23516] == 23516 && 
b[23517] == 23517 && 
b[23518] == 23518 && 
b[23519] == 23519 && 
b[23520] == 23520 && 
b[23521] == 23521 && 
b[23522] == 23522 && 
b[23523] == 23523 && 
b[23524] == 23524 && 
b[23525] == 23525 && 
b[23526] == 23526 && 
b[23527] == 23527 && 
b[23528] == 23528 && 
b[23529] == 23529 && 
b[23530] == 23530 && 
b[23531] == 23531 && 
b[23532] == 23532 && 
b[23533] == 23533 && 
b[23534] == 23534 && 
b[23535] == 23535 && 
b[23536] == 23536 && 
b[23537] == 23537 && 
b[23538] == 23538 && 
b[23539] == 23539 && 
b[23540] == 23540 && 
b[23541] == 23541 && 
b[23542] == 23542 && 
b[23543] == 23543 && 
b[23544] == 23544 && 
b[23545] == 23545 && 
b[23546] == 23546 && 
b[23547] == 23547 && 
b[23548] == 23548 && 
b[23549] == 23549 && 
b[23550] == 23550 && 
b[23551] == 23551 && 
b[23552] == 23552 && 
b[23553] == 23553 && 
b[23554] == 23554 && 
b[23555] == 23555 && 
b[23556] == 23556 && 
b[23557] == 23557 && 
b[23558] == 23558 && 
b[23559] == 23559 && 
b[23560] == 23560 && 
b[23561] == 23561 && 
b[23562] == 23562 && 
b[23563] == 23563 && 
b[23564] == 23564 && 
b[23565] == 23565 && 
b[23566] == 23566 && 
b[23567] == 23567 && 
b[23568] == 23568 && 
b[23569] == 23569 && 
b[23570] == 23570 && 
b[23571] == 23571 && 
b[23572] == 23572 && 
b[23573] == 23573 && 
b[23574] == 23574 && 
b[23575] == 23575 && 
b[23576] == 23576 && 
b[23577] == 23577 && 
b[23578] == 23578 && 
b[23579] == 23579 && 
b[23580] == 23580 && 
b[23581] == 23581 && 
b[23582] == 23582 && 
b[23583] == 23583 && 
b[23584] == 23584 && 
b[23585] == 23585 && 
b[23586] == 23586 && 
b[23587] == 23587 && 
b[23588] == 23588 && 
b[23589] == 23589 && 
b[23590] == 23590 && 
b[23591] == 23591 && 
b[23592] == 23592 && 
b[23593] == 23593 && 
b[23594] == 23594 && 
b[23595] == 23595 && 
b[23596] == 23596 && 
b[23597] == 23597 && 
b[23598] == 23598 && 
b[23599] == 23599 && 
b[23600] == 23600 && 
b[23601] == 23601 && 
b[23602] == 23602 && 
b[23603] == 23603 && 
b[23604] == 23604 && 
b[23605] == 23605 && 
b[23606] == 23606 && 
b[23607] == 23607 && 
b[23608] == 23608 && 
b[23609] == 23609 && 
b[23610] == 23610 && 
b[23611] == 23611 && 
b[23612] == 23612 && 
b[23613] == 23613 && 
b[23614] == 23614 && 
b[23615] == 23615 && 
b[23616] == 23616 && 
b[23617] == 23617 && 
b[23618] == 23618 && 
b[23619] == 23619 && 
b[23620] == 23620 && 
b[23621] == 23621 && 
b[23622] == 23622 && 
b[23623] == 23623 && 
b[23624] == 23624 && 
b[23625] == 23625 && 
b[23626] == 23626 && 
b[23627] == 23627 && 
b[23628] == 23628 && 
b[23629] == 23629 && 
b[23630] == 23630 && 
b[23631] == 23631 && 
b[23632] == 23632 && 
b[23633] == 23633 && 
b[23634] == 23634 && 
b[23635] == 23635 && 
b[23636] == 23636 && 
b[23637] == 23637 && 
b[23638] == 23638 && 
b[23639] == 23639 && 
b[23640] == 23640 && 
b[23641] == 23641 && 
b[23642] == 23642 && 
b[23643] == 23643 && 
b[23644] == 23644 && 
b[23645] == 23645 && 
b[23646] == 23646 && 
b[23647] == 23647 && 
b[23648] == 23648 && 
b[23649] == 23649 && 
b[23650] == 23650 && 
b[23651] == 23651 && 
b[23652] == 23652 && 
b[23653] == 23653 && 
b[23654] == 23654 && 
b[23655] == 23655 && 
b[23656] == 23656 && 
b[23657] == 23657 && 
b[23658] == 23658 && 
b[23659] == 23659 && 
b[23660] == 23660 && 
b[23661] == 23661 && 
b[23662] == 23662 && 
b[23663] == 23663 && 
b[23664] == 23664 && 
b[23665] == 23665 && 
b[23666] == 23666 && 
b[23667] == 23667 && 
b[23668] == 23668 && 
b[23669] == 23669 && 
b[23670] == 23670 && 
b[23671] == 23671 && 
b[23672] == 23672 && 
b[23673] == 23673 && 
b[23674] == 23674 && 
b[23675] == 23675 && 
b[23676] == 23676 && 
b[23677] == 23677 && 
b[23678] == 23678 && 
b[23679] == 23679 && 
b[23680] == 23680 && 
b[23681] == 23681 && 
b[23682] == 23682 && 
b[23683] == 23683 && 
b[23684] == 23684 && 
b[23685] == 23685 && 
b[23686] == 23686 && 
b[23687] == 23687 && 
b[23688] == 23688 && 
b[23689] == 23689 && 
b[23690] == 23690 && 
b[23691] == 23691 && 
b[23692] == 23692 && 
b[23693] == 23693 && 
b[23694] == 23694 && 
b[23695] == 23695 && 
b[23696] == 23696 && 
b[23697] == 23697 && 
b[23698] == 23698 && 
b[23699] == 23699 && 
b[23700] == 23700 && 
b[23701] == 23701 && 
b[23702] == 23702 && 
b[23703] == 23703 && 
b[23704] == 23704 && 
b[23705] == 23705 && 
b[23706] == 23706 && 
b[23707] == 23707 && 
b[23708] == 23708 && 
b[23709] == 23709 && 
b[23710] == 23710 && 
b[23711] == 23711 && 
b[23712] == 23712 && 
b[23713] == 23713 && 
b[23714] == 23714 && 
b[23715] == 23715 && 
b[23716] == 23716 && 
b[23717] == 23717 && 
b[23718] == 23718 && 
b[23719] == 23719 && 
b[23720] == 23720 && 
b[23721] == 23721 && 
b[23722] == 23722 && 
b[23723] == 23723 && 
b[23724] == 23724 && 
b[23725] == 23725 && 
b[23726] == 23726 && 
b[23727] == 23727 && 
b[23728] == 23728 && 
b[23729] == 23729 && 
b[23730] == 23730 && 
b[23731] == 23731 && 
b[23732] == 23732 && 
b[23733] == 23733 && 
b[23734] == 23734 && 
b[23735] == 23735 && 
b[23736] == 23736 && 
b[23737] == 23737 && 
b[23738] == 23738 && 
b[23739] == 23739 && 
b[23740] == 23740 && 
b[23741] == 23741 && 
b[23742] == 23742 && 
b[23743] == 23743 && 
b[23744] == 23744 && 
b[23745] == 23745 && 
b[23746] == 23746 && 
b[23747] == 23747 && 
b[23748] == 23748 && 
b[23749] == 23749 && 
b[23750] == 23750 && 
b[23751] == 23751 && 
b[23752] == 23752 && 
b[23753] == 23753 && 
b[23754] == 23754 && 
b[23755] == 23755 && 
b[23756] == 23756 && 
b[23757] == 23757 && 
b[23758] == 23758 && 
b[23759] == 23759 && 
b[23760] == 23760 && 
b[23761] == 23761 && 
b[23762] == 23762 && 
b[23763] == 23763 && 
b[23764] == 23764 && 
b[23765] == 23765 && 
b[23766] == 23766 && 
b[23767] == 23767 && 
b[23768] == 23768 && 
b[23769] == 23769 && 
b[23770] == 23770 && 
b[23771] == 23771 && 
b[23772] == 23772 && 
b[23773] == 23773 && 
b[23774] == 23774 && 
b[23775] == 23775 && 
b[23776] == 23776 && 
b[23777] == 23777 && 
b[23778] == 23778 && 
b[23779] == 23779 && 
b[23780] == 23780 && 
b[23781] == 23781 && 
b[23782] == 23782 && 
b[23783] == 23783 && 
b[23784] == 23784 && 
b[23785] == 23785 && 
b[23786] == 23786 && 
b[23787] == 23787 && 
b[23788] == 23788 && 
b[23789] == 23789 && 
b[23790] == 23790 && 
b[23791] == 23791 && 
b[23792] == 23792 && 
b[23793] == 23793 && 
b[23794] == 23794 && 
b[23795] == 23795 && 
b[23796] == 23796 && 
b[23797] == 23797 && 
b[23798] == 23798 && 
b[23799] == 23799 && 
b[23800] == 23800 && 
b[23801] == 23801 && 
b[23802] == 23802 && 
b[23803] == 23803 && 
b[23804] == 23804 && 
b[23805] == 23805 && 
b[23806] == 23806 && 
b[23807] == 23807 && 
b[23808] == 23808 && 
b[23809] == 23809 && 
b[23810] == 23810 && 
b[23811] == 23811 && 
b[23812] == 23812 && 
b[23813] == 23813 && 
b[23814] == 23814 && 
b[23815] == 23815 && 
b[23816] == 23816 && 
b[23817] == 23817 && 
b[23818] == 23818 && 
b[23819] == 23819 && 
b[23820] == 23820 && 
b[23821] == 23821 && 
b[23822] == 23822 && 
b[23823] == 23823 && 
b[23824] == 23824 && 
b[23825] == 23825 && 
b[23826] == 23826 && 
b[23827] == 23827 && 
b[23828] == 23828 && 
b[23829] == 23829 && 
b[23830] == 23830 && 
b[23831] == 23831 && 
b[23832] == 23832 && 
b[23833] == 23833 && 
b[23834] == 23834 && 
b[23835] == 23835 && 
b[23836] == 23836 && 
b[23837] == 23837 && 
b[23838] == 23838 && 
b[23839] == 23839 && 
b[23840] == 23840 && 
b[23841] == 23841 && 
b[23842] == 23842 && 
b[23843] == 23843 && 
b[23844] == 23844 && 
b[23845] == 23845 && 
b[23846] == 23846 && 
b[23847] == 23847 && 
b[23848] == 23848 && 
b[23849] == 23849 && 
b[23850] == 23850 && 
b[23851] == 23851 && 
b[23852] == 23852 && 
b[23853] == 23853 && 
b[23854] == 23854 && 
b[23855] == 23855 && 
b[23856] == 23856 && 
b[23857] == 23857 && 
b[23858] == 23858 && 
b[23859] == 23859 && 
b[23860] == 23860 && 
b[23861] == 23861 && 
b[23862] == 23862 && 
b[23863] == 23863 && 
b[23864] == 23864 && 
b[23865] == 23865 && 
b[23866] == 23866 && 
b[23867] == 23867 && 
b[23868] == 23868 && 
b[23869] == 23869 && 
b[23870] == 23870 && 
b[23871] == 23871 && 
b[23872] == 23872 && 
b[23873] == 23873 && 
b[23874] == 23874 && 
b[23875] == 23875 && 
b[23876] == 23876 && 
b[23877] == 23877 && 
b[23878] == 23878 && 
b[23879] == 23879 && 
b[23880] == 23880 && 
b[23881] == 23881 && 
b[23882] == 23882 && 
b[23883] == 23883 && 
b[23884] == 23884 && 
b[23885] == 23885 && 
b[23886] == 23886 && 
b[23887] == 23887 && 
b[23888] == 23888 && 
b[23889] == 23889 && 
b[23890] == 23890 && 
b[23891] == 23891 && 
b[23892] == 23892 && 
b[23893] == 23893 && 
b[23894] == 23894 && 
b[23895] == 23895 && 
b[23896] == 23896 && 
b[23897] == 23897 && 
b[23898] == 23898 && 
b[23899] == 23899 && 
b[23900] == 23900 && 
b[23901] == 23901 && 
b[23902] == 23902 && 
b[23903] == 23903 && 
b[23904] == 23904 && 
b[23905] == 23905 && 
b[23906] == 23906 && 
b[23907] == 23907 && 
b[23908] == 23908 && 
b[23909] == 23909 && 
b[23910] == 23910 && 
b[23911] == 23911 && 
b[23912] == 23912 && 
b[23913] == 23913 && 
b[23914] == 23914 && 
b[23915] == 23915 && 
b[23916] == 23916 && 
b[23917] == 23917 && 
b[23918] == 23918 && 
b[23919] == 23919 && 
b[23920] == 23920 && 
b[23921] == 23921 && 
b[23922] == 23922 && 
b[23923] == 23923 && 
b[23924] == 23924 && 
b[23925] == 23925 && 
b[23926] == 23926 && 
b[23927] == 23927 && 
b[23928] == 23928 && 
b[23929] == 23929 && 
b[23930] == 23930 && 
b[23931] == 23931 && 
b[23932] == 23932 && 
b[23933] == 23933 && 
b[23934] == 23934 && 
b[23935] == 23935 && 
b[23936] == 23936 && 
b[23937] == 23937 && 
b[23938] == 23938 && 
b[23939] == 23939 && 
b[23940] == 23940 && 
b[23941] == 23941 && 
b[23942] == 23942 && 
b[23943] == 23943 && 
b[23944] == 23944 && 
b[23945] == 23945 && 
b[23946] == 23946 && 
b[23947] == 23947 && 
b[23948] == 23948 && 
b[23949] == 23949 && 
b[23950] == 23950 && 
b[23951] == 23951 && 
b[23952] == 23952 && 
b[23953] == 23953 && 
b[23954] == 23954 && 
b[23955] == 23955 && 
b[23956] == 23956 && 
b[23957] == 23957 && 
b[23958] == 23958 && 
b[23959] == 23959 && 
b[23960] == 23960 && 
b[23961] == 23961 && 
b[23962] == 23962 && 
b[23963] == 23963 && 
b[23964] == 23964 && 
b[23965] == 23965 && 
b[23966] == 23966 && 
b[23967] == 23967 && 
b[23968] == 23968 && 
b[23969] == 23969 && 
b[23970] == 23970 && 
b[23971] == 23971 && 
b[23972] == 23972 && 
b[23973] == 23973 && 
b[23974] == 23974 && 
b[23975] == 23975 && 
b[23976] == 23976 && 
b[23977] == 23977 && 
b[23978] == 23978 && 
b[23979] == 23979 && 
b[23980] == 23980 && 
b[23981] == 23981 && 
b[23982] == 23982 && 
b[23983] == 23983 && 
b[23984] == 23984 && 
b[23985] == 23985 && 
b[23986] == 23986 && 
b[23987] == 23987 && 
b[23988] == 23988 && 
b[23989] == 23989 && 
b[23990] == 23990 && 
b[23991] == 23991 && 
b[23992] == 23992 && 
b[23993] == 23993 && 
b[23994] == 23994 && 
b[23995] == 23995 && 
b[23996] == 23996 && 
b[23997] == 23997 && 
b[23998] == 23998 && 
b[23999] == 23999 && 
b[24000] == 24000 && 
b[24001] == 24001 && 
b[24002] == 24002 && 
b[24003] == 24003 && 
b[24004] == 24004 && 
b[24005] == 24005 && 
b[24006] == 24006 && 
b[24007] == 24007 && 
b[24008] == 24008 && 
b[24009] == 24009 && 
b[24010] == 24010 && 
b[24011] == 24011 && 
b[24012] == 24012 && 
b[24013] == 24013 && 
b[24014] == 24014 && 
b[24015] == 24015 && 
b[24016] == 24016 && 
b[24017] == 24017 && 
b[24018] == 24018 && 
b[24019] == 24019 && 
b[24020] == 24020 && 
b[24021] == 24021 && 
b[24022] == 24022 && 
b[24023] == 24023 && 
b[24024] == 24024 && 
b[24025] == 24025 && 
b[24026] == 24026 && 
b[24027] == 24027 && 
b[24028] == 24028 && 
b[24029] == 24029 && 
b[24030] == 24030 && 
b[24031] == 24031 && 
b[24032] == 24032 && 
b[24033] == 24033 && 
b[24034] == 24034 && 
b[24035] == 24035 && 
b[24036] == 24036 && 
b[24037] == 24037 && 
b[24038] == 24038 && 
b[24039] == 24039 && 
b[24040] == 24040 && 
b[24041] == 24041 && 
b[24042] == 24042 && 
b[24043] == 24043 && 
b[24044] == 24044 && 
b[24045] == 24045 && 
b[24046] == 24046 && 
b[24047] == 24047 && 
b[24048] == 24048 && 
b[24049] == 24049 && 
b[24050] == 24050 && 
b[24051] == 24051 && 
b[24052] == 24052 && 
b[24053] == 24053 && 
b[24054] == 24054 && 
b[24055] == 24055 && 
b[24056] == 24056 && 
b[24057] == 24057 && 
b[24058] == 24058 && 
b[24059] == 24059 && 
b[24060] == 24060 && 
b[24061] == 24061 && 
b[24062] == 24062 && 
b[24063] == 24063 && 
b[24064] == 24064 && 
b[24065] == 24065 && 
b[24066] == 24066 && 
b[24067] == 24067 && 
b[24068] == 24068 && 
b[24069] == 24069 && 
b[24070] == 24070 && 
b[24071] == 24071 && 
b[24072] == 24072 && 
b[24073] == 24073 && 
b[24074] == 24074 && 
b[24075] == 24075 && 
b[24076] == 24076 && 
b[24077] == 24077 && 
b[24078] == 24078 && 
b[24079] == 24079 && 
b[24080] == 24080 && 
b[24081] == 24081 && 
b[24082] == 24082 && 
b[24083] == 24083 && 
b[24084] == 24084 && 
b[24085] == 24085 && 
b[24086] == 24086 && 
b[24087] == 24087 && 
b[24088] == 24088 && 
b[24089] == 24089 && 
b[24090] == 24090 && 
b[24091] == 24091 && 
b[24092] == 24092 && 
b[24093] == 24093 && 
b[24094] == 24094 && 
b[24095] == 24095 && 
b[24096] == 24096 && 
b[24097] == 24097 && 
b[24098] == 24098 && 
b[24099] == 24099 && 
b[24100] == 24100 && 
b[24101] == 24101 && 
b[24102] == 24102 && 
b[24103] == 24103 && 
b[24104] == 24104 && 
b[24105] == 24105 && 
b[24106] == 24106 && 
b[24107] == 24107 && 
b[24108] == 24108 && 
b[24109] == 24109 && 
b[24110] == 24110 && 
b[24111] == 24111 && 
b[24112] == 24112 && 
b[24113] == 24113 && 
b[24114] == 24114 && 
b[24115] == 24115 && 
b[24116] == 24116 && 
b[24117] == 24117 && 
b[24118] == 24118 && 
b[24119] == 24119 && 
b[24120] == 24120 && 
b[24121] == 24121 && 
b[24122] == 24122 && 
b[24123] == 24123 && 
b[24124] == 24124 && 
b[24125] == 24125 && 
b[24126] == 24126 && 
b[24127] == 24127 && 
b[24128] == 24128 && 
b[24129] == 24129 && 
b[24130] == 24130 && 
b[24131] == 24131 && 
b[24132] == 24132 && 
b[24133] == 24133 && 
b[24134] == 24134 && 
b[24135] == 24135 && 
b[24136] == 24136 && 
b[24137] == 24137 && 
b[24138] == 24138 && 
b[24139] == 24139 && 
b[24140] == 24140 && 
b[24141] == 24141 && 
b[24142] == 24142 && 
b[24143] == 24143 && 
b[24144] == 24144 && 
b[24145] == 24145 && 
b[24146] == 24146 && 
b[24147] == 24147 && 
b[24148] == 24148 && 
b[24149] == 24149 && 
b[24150] == 24150 && 
b[24151] == 24151 && 
b[24152] == 24152 && 
b[24153] == 24153 && 
b[24154] == 24154 && 
b[24155] == 24155 && 
b[24156] == 24156 && 
b[24157] == 24157 && 
b[24158] == 24158 && 
b[24159] == 24159 && 
b[24160] == 24160 && 
b[24161] == 24161 && 
b[24162] == 24162 && 
b[24163] == 24163 && 
b[24164] == 24164 && 
b[24165] == 24165 && 
b[24166] == 24166 && 
b[24167] == 24167 && 
b[24168] == 24168 && 
b[24169] == 24169 && 
b[24170] == 24170 && 
b[24171] == 24171 && 
b[24172] == 24172 && 
b[24173] == 24173 && 
b[24174] == 24174 && 
b[24175] == 24175 && 
b[24176] == 24176 && 
b[24177] == 24177 && 
b[24178] == 24178 && 
b[24179] == 24179 && 
b[24180] == 24180 && 
b[24181] == 24181 && 
b[24182] == 24182 && 
b[24183] == 24183 && 
b[24184] == 24184 && 
b[24185] == 24185 && 
b[24186] == 24186 && 
b[24187] == 24187 && 
b[24188] == 24188 && 
b[24189] == 24189 && 
b[24190] == 24190 && 
b[24191] == 24191 && 
b[24192] == 24192 && 
b[24193] == 24193 && 
b[24194] == 24194 && 
b[24195] == 24195 && 
b[24196] == 24196 && 
b[24197] == 24197 && 
b[24198] == 24198 && 
b[24199] == 24199 && 
b[24200] == 24200 && 
b[24201] == 24201 && 
b[24202] == 24202 && 
b[24203] == 24203 && 
b[24204] == 24204 && 
b[24205] == 24205 && 
b[24206] == 24206 && 
b[24207] == 24207 && 
b[24208] == 24208 && 
b[24209] == 24209 && 
b[24210] == 24210 && 
b[24211] == 24211 && 
b[24212] == 24212 && 
b[24213] == 24213 && 
b[24214] == 24214 && 
b[24215] == 24215 && 
b[24216] == 24216 && 
b[24217] == 24217 && 
b[24218] == 24218 && 
b[24219] == 24219 && 
b[24220] == 24220 && 
b[24221] == 24221 && 
b[24222] == 24222 && 
b[24223] == 24223 && 
b[24224] == 24224 && 
b[24225] == 24225 && 
b[24226] == 24226 && 
b[24227] == 24227 && 
b[24228] == 24228 && 
b[24229] == 24229 && 
b[24230] == 24230 && 
b[24231] == 24231 && 
b[24232] == 24232 && 
b[24233] == 24233 && 
b[24234] == 24234 && 
b[24235] == 24235 && 
b[24236] == 24236 && 
b[24237] == 24237 && 
b[24238] == 24238 && 
b[24239] == 24239 && 
b[24240] == 24240 && 
b[24241] == 24241 && 
b[24242] == 24242 && 
b[24243] == 24243 && 
b[24244] == 24244 && 
b[24245] == 24245 && 
b[24246] == 24246 && 
b[24247] == 24247 && 
b[24248] == 24248 && 
b[24249] == 24249 && 
b[24250] == 24250 && 
b[24251] == 24251 && 
b[24252] == 24252 && 
b[24253] == 24253 && 
b[24254] == 24254 && 
b[24255] == 24255 && 
b[24256] == 24256 && 
b[24257] == 24257 && 
b[24258] == 24258 && 
b[24259] == 24259 && 
b[24260] == 24260 && 
b[24261] == 24261 && 
b[24262] == 24262 && 
b[24263] == 24263 && 
b[24264] == 24264 && 
b[24265] == 24265 && 
b[24266] == 24266 && 
b[24267] == 24267 && 
b[24268] == 24268 && 
b[24269] == 24269 && 
b[24270] == 24270 && 
b[24271] == 24271 && 
b[24272] == 24272 && 
b[24273] == 24273 && 
b[24274] == 24274 && 
b[24275] == 24275 && 
b[24276] == 24276 && 
b[24277] == 24277 && 
b[24278] == 24278 && 
b[24279] == 24279 && 
b[24280] == 24280 && 
b[24281] == 24281 && 
b[24282] == 24282 && 
b[24283] == 24283 && 
b[24284] == 24284 && 
b[24285] == 24285 && 
b[24286] == 24286 && 
b[24287] == 24287 && 
b[24288] == 24288 && 
b[24289] == 24289 && 
b[24290] == 24290 && 
b[24291] == 24291 && 
b[24292] == 24292 && 
b[24293] == 24293 && 
b[24294] == 24294 && 
b[24295] == 24295 && 
b[24296] == 24296 && 
b[24297] == 24297 && 
b[24298] == 24298 && 
b[24299] == 24299 && 
b[24300] == 24300 && 
b[24301] == 24301 && 
b[24302] == 24302 && 
b[24303] == 24303 && 
b[24304] == 24304 && 
b[24305] == 24305 && 
b[24306] == 24306 && 
b[24307] == 24307 && 
b[24308] == 24308 && 
b[24309] == 24309 && 
b[24310] == 24310 && 
b[24311] == 24311 && 
b[24312] == 24312 && 
b[24313] == 24313 && 
b[24314] == 24314 && 
b[24315] == 24315 && 
b[24316] == 24316 && 
b[24317] == 24317 && 
b[24318] == 24318 && 
b[24319] == 24319 && 
b[24320] == 24320 && 
b[24321] == 24321 && 
b[24322] == 24322 && 
b[24323] == 24323 && 
b[24324] == 24324 && 
b[24325] == 24325 && 
b[24326] == 24326 && 
b[24327] == 24327 && 
b[24328] == 24328 && 
b[24329] == 24329 && 
b[24330] == 24330 && 
b[24331] == 24331 && 
b[24332] == 24332 && 
b[24333] == 24333 && 
b[24334] == 24334 && 
b[24335] == 24335 && 
b[24336] == 24336 && 
b[24337] == 24337 && 
b[24338] == 24338 && 
b[24339] == 24339 && 
b[24340] == 24340 && 
b[24341] == 24341 && 
b[24342] == 24342 && 
b[24343] == 24343 && 
b[24344] == 24344 && 
b[24345] == 24345 && 
b[24346] == 24346 && 
b[24347] == 24347 && 
b[24348] == 24348 && 
b[24349] == 24349 && 
b[24350] == 24350 && 
b[24351] == 24351 && 
b[24352] == 24352 && 
b[24353] == 24353 && 
b[24354] == 24354 && 
b[24355] == 24355 && 
b[24356] == 24356 && 
b[24357] == 24357 && 
b[24358] == 24358 && 
b[24359] == 24359 && 
b[24360] == 24360 && 
b[24361] == 24361 && 
b[24362] == 24362 && 
b[24363] == 24363 && 
b[24364] == 24364 && 
b[24365] == 24365 && 
b[24366] == 24366 && 
b[24367] == 24367 && 
b[24368] == 24368 && 
b[24369] == 24369 && 
b[24370] == 24370 && 
b[24371] == 24371 && 
b[24372] == 24372 && 
b[24373] == 24373 && 
b[24374] == 24374 && 
b[24375] == 24375 && 
b[24376] == 24376 && 
b[24377] == 24377 && 
b[24378] == 24378 && 
b[24379] == 24379 && 
b[24380] == 24380 && 
b[24381] == 24381 && 
b[24382] == 24382 && 
b[24383] == 24383 && 
b[24384] == 24384 && 
b[24385] == 24385 && 
b[24386] == 24386 && 
b[24387] == 24387 && 
b[24388] == 24388 && 
b[24389] == 24389 && 
b[24390] == 24390 && 
b[24391] == 24391 && 
b[24392] == 24392 && 
b[24393] == 24393 && 
b[24394] == 24394 && 
b[24395] == 24395 && 
b[24396] == 24396 && 
b[24397] == 24397 && 
b[24398] == 24398 && 
b[24399] == 24399 && 
b[24400] == 24400 && 
b[24401] == 24401 && 
b[24402] == 24402 && 
b[24403] == 24403 && 
b[24404] == 24404 && 
b[24405] == 24405 && 
b[24406] == 24406 && 
b[24407] == 24407 && 
b[24408] == 24408 && 
b[24409] == 24409 && 
b[24410] == 24410 && 
b[24411] == 24411 && 
b[24412] == 24412 && 
b[24413] == 24413 && 
b[24414] == 24414 && 
b[24415] == 24415 && 
b[24416] == 24416 && 
b[24417] == 24417 && 
b[24418] == 24418 && 
b[24419] == 24419 && 
b[24420] == 24420 && 
b[24421] == 24421 && 
b[24422] == 24422 && 
b[24423] == 24423 && 
b[24424] == 24424 && 
b[24425] == 24425 && 
b[24426] == 24426 && 
b[24427] == 24427 && 
b[24428] == 24428 && 
b[24429] == 24429 && 
b[24430] == 24430 && 
b[24431] == 24431 && 
b[24432] == 24432 && 
b[24433] == 24433 && 
b[24434] == 24434 && 
b[24435] == 24435 && 
b[24436] == 24436 && 
b[24437] == 24437 && 
b[24438] == 24438 && 
b[24439] == 24439 && 
b[24440] == 24440 && 
b[24441] == 24441 && 
b[24442] == 24442 && 
b[24443] == 24443 && 
b[24444] == 24444 && 
b[24445] == 24445 && 
b[24446] == 24446 && 
b[24447] == 24447 && 
b[24448] == 24448 && 
b[24449] == 24449 && 
b[24450] == 24450 && 
b[24451] == 24451 && 
b[24452] == 24452 && 
b[24453] == 24453 && 
b[24454] == 24454 && 
b[24455] == 24455 && 
b[24456] == 24456 && 
b[24457] == 24457 && 
b[24458] == 24458 && 
b[24459] == 24459 && 
b[24460] == 24460 && 
b[24461] == 24461 && 
b[24462] == 24462 && 
b[24463] == 24463 && 
b[24464] == 24464 && 
b[24465] == 24465 && 
b[24466] == 24466 && 
b[24467] == 24467 && 
b[24468] == 24468 && 
b[24469] == 24469 && 
b[24470] == 24470 && 
b[24471] == 24471 && 
b[24472] == 24472 && 
b[24473] == 24473 && 
b[24474] == 24474 && 
b[24475] == 24475 && 
b[24476] == 24476 && 
b[24477] == 24477 && 
b[24478] == 24478 && 
b[24479] == 24479 && 
b[24480] == 24480 && 
b[24481] == 24481 && 
b[24482] == 24482 && 
b[24483] == 24483 && 
b[24484] == 24484 && 
b[24485] == 24485 && 
b[24486] == 24486 && 
b[24487] == 24487 && 
b[24488] == 24488 && 
b[24489] == 24489 && 
b[24490] == 24490 && 
b[24491] == 24491 && 
b[24492] == 24492 && 
b[24493] == 24493 && 
b[24494] == 24494 && 
b[24495] == 24495 && 
b[24496] == 24496 && 
b[24497] == 24497 && 
b[24498] == 24498 && 
b[24499] == 24499 && 
b[24500] == 24500 && 
b[24501] == 24501 && 
b[24502] == 24502 && 
b[24503] == 24503 && 
b[24504] == 24504 && 
b[24505] == 24505 && 
b[24506] == 24506 && 
b[24507] == 24507 && 
b[24508] == 24508 && 
b[24509] == 24509 && 
b[24510] == 24510 && 
b[24511] == 24511 && 
b[24512] == 24512 && 
b[24513] == 24513 && 
b[24514] == 24514 && 
b[24515] == 24515 && 
b[24516] == 24516 && 
b[24517] == 24517 && 
b[24518] == 24518 && 
b[24519] == 24519 && 
b[24520] == 24520 && 
b[24521] == 24521 && 
b[24522] == 24522 && 
b[24523] == 24523 && 
b[24524] == 24524 && 
b[24525] == 24525 && 
b[24526] == 24526 && 
b[24527] == 24527 && 
b[24528] == 24528 && 
b[24529] == 24529 && 
b[24530] == 24530 && 
b[24531] == 24531 && 
b[24532] == 24532 && 
b[24533] == 24533 && 
b[24534] == 24534 && 
b[24535] == 24535 && 
b[24536] == 24536 && 
b[24537] == 24537 && 
b[24538] == 24538 && 
b[24539] == 24539 && 
b[24540] == 24540 && 
b[24541] == 24541 && 
b[24542] == 24542 && 
b[24543] == 24543 && 
b[24544] == 24544 && 
b[24545] == 24545 && 
b[24546] == 24546 && 
b[24547] == 24547 && 
b[24548] == 24548 && 
b[24549] == 24549 && 
b[24550] == 24550 && 
b[24551] == 24551 && 
b[24552] == 24552 && 
b[24553] == 24553 && 
b[24554] == 24554 && 
b[24555] == 24555 && 
b[24556] == 24556 && 
b[24557] == 24557 && 
b[24558] == 24558 && 
b[24559] == 24559 && 
b[24560] == 24560 && 
b[24561] == 24561 && 
b[24562] == 24562 && 
b[24563] == 24563 && 
b[24564] == 24564 && 
b[24565] == 24565 && 
b[24566] == 24566 && 
b[24567] == 24567 && 
b[24568] == 24568 && 
b[24569] == 24569 && 
b[24570] == 24570 && 
b[24571] == 24571 && 
b[24572] == 24572 && 
b[24573] == 24573 && 
b[24574] == 24574 && 
b[24575] == 24575 && 
b[24576] == 24576 && 
b[24577] == 24577 && 
b[24578] == 24578 && 
b[24579] == 24579 && 
b[24580] == 24580 && 
b[24581] == 24581 && 
b[24582] == 24582 && 
b[24583] == 24583 && 
b[24584] == 24584 && 
b[24585] == 24585 && 
b[24586] == 24586 && 
b[24587] == 24587 && 
b[24588] == 24588 && 
b[24589] == 24589 && 
b[24590] == 24590 && 
b[24591] == 24591 && 
b[24592] == 24592 && 
b[24593] == 24593 && 
b[24594] == 24594 && 
b[24595] == 24595 && 
b[24596] == 24596 && 
b[24597] == 24597 && 
b[24598] == 24598 && 
b[24599] == 24599 && 
b[24600] == 24600 && 
b[24601] == 24601 && 
b[24602] == 24602 && 
b[24603] == 24603 && 
b[24604] == 24604 && 
b[24605] == 24605 && 
b[24606] == 24606 && 
b[24607] == 24607 && 
b[24608] == 24608 && 
b[24609] == 24609 && 
b[24610] == 24610 && 
b[24611] == 24611 && 
b[24612] == 24612 && 
b[24613] == 24613 && 
b[24614] == 24614 && 
b[24615] == 24615 && 
b[24616] == 24616 && 
b[24617] == 24617 && 
b[24618] == 24618 && 
b[24619] == 24619 && 
b[24620] == 24620 && 
b[24621] == 24621 && 
b[24622] == 24622 && 
b[24623] == 24623 && 
b[24624] == 24624 && 
b[24625] == 24625 && 
b[24626] == 24626 && 
b[24627] == 24627 && 
b[24628] == 24628 && 
b[24629] == 24629 && 
b[24630] == 24630 && 
b[24631] == 24631 && 
b[24632] == 24632 && 
b[24633] == 24633 && 
b[24634] == 24634 && 
b[24635] == 24635 && 
b[24636] == 24636 && 
b[24637] == 24637 && 
b[24638] == 24638 && 
b[24639] == 24639 && 
b[24640] == 24640 && 
b[24641] == 24641 && 
b[24642] == 24642 && 
b[24643] == 24643 && 
b[24644] == 24644 && 
b[24645] == 24645 && 
b[24646] == 24646 && 
b[24647] == 24647 && 
b[24648] == 24648 && 
b[24649] == 24649 && 
b[24650] == 24650 && 
b[24651] == 24651 && 
b[24652] == 24652 && 
b[24653] == 24653 && 
b[24654] == 24654 && 
b[24655] == 24655 && 
b[24656] == 24656 && 
b[24657] == 24657 && 
b[24658] == 24658 && 
b[24659] == 24659 && 
b[24660] == 24660 && 
b[24661] == 24661 && 
b[24662] == 24662 && 
b[24663] == 24663 && 
b[24664] == 24664 && 
b[24665] == 24665 && 
b[24666] == 24666 && 
b[24667] == 24667 && 
b[24668] == 24668 && 
b[24669] == 24669 && 
b[24670] == 24670 && 
b[24671] == 24671 && 
b[24672] == 24672 && 
b[24673] == 24673 && 
b[24674] == 24674 && 
b[24675] == 24675 && 
b[24676] == 24676 && 
b[24677] == 24677 && 
b[24678] == 24678 && 
b[24679] == 24679 && 
b[24680] == 24680 && 
b[24681] == 24681 && 
b[24682] == 24682 && 
b[24683] == 24683 && 
b[24684] == 24684 && 
b[24685] == 24685 && 
b[24686] == 24686 && 
b[24687] == 24687 && 
b[24688] == 24688 && 
b[24689] == 24689 && 
b[24690] == 24690 && 
b[24691] == 24691 && 
b[24692] == 24692 && 
b[24693] == 24693 && 
b[24694] == 24694 && 
b[24695] == 24695 && 
b[24696] == 24696 && 
b[24697] == 24697 && 
b[24698] == 24698 && 
b[24699] == 24699 && 
b[24700] == 24700 && 
b[24701] == 24701 && 
b[24702] == 24702 && 
b[24703] == 24703 && 
b[24704] == 24704 && 
b[24705] == 24705 && 
b[24706] == 24706 && 
b[24707] == 24707 && 
b[24708] == 24708 && 
b[24709] == 24709 && 
b[24710] == 24710 && 
b[24711] == 24711 && 
b[24712] == 24712 && 
b[24713] == 24713 && 
b[24714] == 24714 && 
b[24715] == 24715 && 
b[24716] == 24716 && 
b[24717] == 24717 && 
b[24718] == 24718 && 
b[24719] == 24719 && 
b[24720] == 24720 && 
b[24721] == 24721 && 
b[24722] == 24722 && 
b[24723] == 24723 && 
b[24724] == 24724 && 
b[24725] == 24725 && 
b[24726] == 24726 && 
b[24727] == 24727 && 
b[24728] == 24728 && 
b[24729] == 24729 && 
b[24730] == 24730 && 
b[24731] == 24731 && 
b[24732] == 24732 && 
b[24733] == 24733 && 
b[24734] == 24734 && 
b[24735] == 24735 && 
b[24736] == 24736 && 
b[24737] == 24737 && 
b[24738] == 24738 && 
b[24739] == 24739 && 
b[24740] == 24740 && 
b[24741] == 24741 && 
b[24742] == 24742 && 
b[24743] == 24743 && 
b[24744] == 24744 && 
b[24745] == 24745 && 
b[24746] == 24746 && 
b[24747] == 24747 && 
b[24748] == 24748 && 
b[24749] == 24749 && 
b[24750] == 24750 && 
b[24751] == 24751 && 
b[24752] == 24752 && 
b[24753] == 24753 && 
b[24754] == 24754 && 
b[24755] == 24755 && 
b[24756] == 24756 && 
b[24757] == 24757 && 
b[24758] == 24758 && 
b[24759] == 24759 && 
b[24760] == 24760 && 
b[24761] == 24761 && 
b[24762] == 24762 && 
b[24763] == 24763 && 
b[24764] == 24764 && 
b[24765] == 24765 && 
b[24766] == 24766 && 
b[24767] == 24767 && 
b[24768] == 24768 && 
b[24769] == 24769 && 
b[24770] == 24770 && 
b[24771] == 24771 && 
b[24772] == 24772 && 
b[24773] == 24773 && 
b[24774] == 24774 && 
b[24775] == 24775 && 
b[24776] == 24776 && 
b[24777] == 24777 && 
b[24778] == 24778 && 
b[24779] == 24779 && 
b[24780] == 24780 && 
b[24781] == 24781 && 
b[24782] == 24782 && 
b[24783] == 24783 && 
b[24784] == 24784 && 
b[24785] == 24785 && 
b[24786] == 24786 && 
b[24787] == 24787 && 
b[24788] == 24788 && 
b[24789] == 24789 && 
b[24790] == 24790 && 
b[24791] == 24791 && 
b[24792] == 24792 && 
b[24793] == 24793 && 
b[24794] == 24794 && 
b[24795] == 24795 && 
b[24796] == 24796 && 
b[24797] == 24797 && 
b[24798] == 24798 && 
b[24799] == 24799 && 
b[24800] == 24800 && 
b[24801] == 24801 && 
b[24802] == 24802 && 
b[24803] == 24803 && 
b[24804] == 24804 && 
b[24805] == 24805 && 
b[24806] == 24806 && 
b[24807] == 24807 && 
b[24808] == 24808 && 
b[24809] == 24809 && 
b[24810] == 24810 && 
b[24811] == 24811 && 
b[24812] == 24812 && 
b[24813] == 24813 && 
b[24814] == 24814 && 
b[24815] == 24815 && 
b[24816] == 24816 && 
b[24817] == 24817 && 
b[24818] == 24818 && 
b[24819] == 24819 && 
b[24820] == 24820 && 
b[24821] == 24821 && 
b[24822] == 24822 && 
b[24823] == 24823 && 
b[24824] == 24824 && 
b[24825] == 24825 && 
b[24826] == 24826 && 
b[24827] == 24827 && 
b[24828] == 24828 && 
b[24829] == 24829 && 
b[24830] == 24830 && 
b[24831] == 24831 && 
b[24832] == 24832 && 
b[24833] == 24833 && 
b[24834] == 24834 && 
b[24835] == 24835 && 
b[24836] == 24836 && 
b[24837] == 24837 && 
b[24838] == 24838 && 
b[24839] == 24839 && 
b[24840] == 24840 && 
b[24841] == 24841 && 
b[24842] == 24842 && 
b[24843] == 24843 && 
b[24844] == 24844 && 
b[24845] == 24845 && 
b[24846] == 24846 && 
b[24847] == 24847 && 
b[24848] == 24848 && 
b[24849] == 24849 && 
b[24850] == 24850 && 
b[24851] == 24851 && 
b[24852] == 24852 && 
b[24853] == 24853 && 
b[24854] == 24854 && 
b[24855] == 24855 && 
b[24856] == 24856 && 
b[24857] == 24857 && 
b[24858] == 24858 && 
b[24859] == 24859 && 
b[24860] == 24860 && 
b[24861] == 24861 && 
b[24862] == 24862 && 
b[24863] == 24863 && 
b[24864] == 24864 && 
b[24865] == 24865 && 
b[24866] == 24866 && 
b[24867] == 24867 && 
b[24868] == 24868 && 
b[24869] == 24869 && 
b[24870] == 24870 && 
b[24871] == 24871 && 
b[24872] == 24872 && 
b[24873] == 24873 && 
b[24874] == 24874 && 
b[24875] == 24875 && 
b[24876] == 24876 && 
b[24877] == 24877 && 
b[24878] == 24878 && 
b[24879] == 24879 && 
b[24880] == 24880 && 
b[24881] == 24881 && 
b[24882] == 24882 && 
b[24883] == 24883 && 
b[24884] == 24884 && 
b[24885] == 24885 && 
b[24886] == 24886 && 
b[24887] == 24887 && 
b[24888] == 24888 && 
b[24889] == 24889 && 
b[24890] == 24890 && 
b[24891] == 24891 && 
b[24892] == 24892 && 
b[24893] == 24893 && 
b[24894] == 24894 && 
b[24895] == 24895 && 
b[24896] == 24896 && 
b[24897] == 24897 && 
b[24898] == 24898 && 
b[24899] == 24899 && 
b[24900] == 24900 && 
b[24901] == 24901 && 
b[24902] == 24902 && 
b[24903] == 24903 && 
b[24904] == 24904 && 
b[24905] == 24905 && 
b[24906] == 24906 && 
b[24907] == 24907 && 
b[24908] == 24908 && 
b[24909] == 24909 && 
b[24910] == 24910 && 
b[24911] == 24911 && 
b[24912] == 24912 && 
b[24913] == 24913 && 
b[24914] == 24914 && 
b[24915] == 24915 && 
b[24916] == 24916 && 
b[24917] == 24917 && 
b[24918] == 24918 && 
b[24919] == 24919 && 
b[24920] == 24920 && 
b[24921] == 24921 && 
b[24922] == 24922 && 
b[24923] == 24923 && 
b[24924] == 24924 && 
b[24925] == 24925 && 
b[24926] == 24926 && 
b[24927] == 24927 && 
b[24928] == 24928 && 
b[24929] == 24929 && 
b[24930] == 24930 && 
b[24931] == 24931 && 
b[24932] == 24932 && 
b[24933] == 24933 && 
b[24934] == 24934 && 
b[24935] == 24935 && 
b[24936] == 24936 && 
b[24937] == 24937 && 
b[24938] == 24938 && 
b[24939] == 24939 && 
b[24940] == 24940 && 
b[24941] == 24941 && 
b[24942] == 24942 && 
b[24943] == 24943 && 
b[24944] == 24944 && 
b[24945] == 24945 && 
b[24946] == 24946 && 
b[24947] == 24947 && 
b[24948] == 24948 && 
b[24949] == 24949 && 
b[24950] == 24950 && 
b[24951] == 24951 && 
b[24952] == 24952 && 
b[24953] == 24953 && 
b[24954] == 24954 && 
b[24955] == 24955 && 
b[24956] == 24956 && 
b[24957] == 24957 && 
b[24958] == 24958 && 
b[24959] == 24959 && 
b[24960] == 24960 && 
b[24961] == 24961 && 
b[24962] == 24962 && 
b[24963] == 24963 && 
b[24964] == 24964 && 
b[24965] == 24965 && 
b[24966] == 24966 && 
b[24967] == 24967 && 
b[24968] == 24968 && 
b[24969] == 24969 && 
b[24970] == 24970 && 
b[24971] == 24971 && 
b[24972] == 24972 && 
b[24973] == 24973 && 
b[24974] == 24974 && 
b[24975] == 24975 && 
b[24976] == 24976 && 
b[24977] == 24977 && 
b[24978] == 24978 && 
b[24979] == 24979 && 
b[24980] == 24980 && 
b[24981] == 24981 && 
b[24982] == 24982 && 
b[24983] == 24983 && 
b[24984] == 24984 && 
b[24985] == 24985 && 
b[24986] == 24986 && 
b[24987] == 24987 && 
b[24988] == 24988 && 
b[24989] == 24989 && 
b[24990] == 24990 && 
b[24991] == 24991 && 
b[24992] == 24992 && 
b[24993] == 24993 && 
b[24994] == 24994 && 
b[24995] == 24995 && 
b[24996] == 24996 && 
b[24997] == 24997 && 
b[24998] == 24998 && 
b[24999] == 24999 && 
b[25000] == 25000 && 
b[25001] == 25001 && 
b[25002] == 25002 && 
b[25003] == 25003 && 
b[25004] == 25004 && 
b[25005] == 25005 && 
b[25006] == 25006 && 
b[25007] == 25007 && 
b[25008] == 25008 && 
b[25009] == 25009 && 
b[25010] == 25010 && 
b[25011] == 25011 && 
b[25012] == 25012 && 
b[25013] == 25013 && 
b[25014] == 25014 && 
b[25015] == 25015 && 
b[25016] == 25016 && 
b[25017] == 25017 && 
b[25018] == 25018 && 
b[25019] == 25019 && 
b[25020] == 25020 && 
b[25021] == 25021 && 
b[25022] == 25022 && 
b[25023] == 25023 && 
b[25024] == 25024 && 
b[25025] == 25025 && 
b[25026] == 25026 && 
b[25027] == 25027 && 
b[25028] == 25028 && 
b[25029] == 25029 && 
b[25030] == 25030 && 
b[25031] == 25031 && 
b[25032] == 25032 && 
b[25033] == 25033 && 
b[25034] == 25034 && 
b[25035] == 25035 && 
b[25036] == 25036 && 
b[25037] == 25037 && 
b[25038] == 25038 && 
b[25039] == 25039 && 
b[25040] == 25040 && 
b[25041] == 25041 && 
b[25042] == 25042 && 
b[25043] == 25043 && 
b[25044] == 25044 && 
b[25045] == 25045 && 
b[25046] == 25046 && 
b[25047] == 25047 && 
b[25048] == 25048 && 
b[25049] == 25049 && 
b[25050] == 25050 && 
b[25051] == 25051 && 
b[25052] == 25052 && 
b[25053] == 25053 && 
b[25054] == 25054 && 
b[25055] == 25055 && 
b[25056] == 25056 && 
b[25057] == 25057 && 
b[25058] == 25058 && 
b[25059] == 25059 && 
b[25060] == 25060 && 
b[25061] == 25061 && 
b[25062] == 25062 && 
b[25063] == 25063 && 
b[25064] == 25064 && 
b[25065] == 25065 && 
b[25066] == 25066 && 
b[25067] == 25067 && 
b[25068] == 25068 && 
b[25069] == 25069 && 
b[25070] == 25070 && 
b[25071] == 25071 && 
b[25072] == 25072 && 
b[25073] == 25073 && 
b[25074] == 25074 && 
b[25075] == 25075 && 
b[25076] == 25076 && 
b[25077] == 25077 && 
b[25078] == 25078 && 
b[25079] == 25079 && 
b[25080] == 25080 && 
b[25081] == 25081 && 
b[25082] == 25082 && 
b[25083] == 25083 && 
b[25084] == 25084 && 
b[25085] == 25085 && 
b[25086] == 25086 && 
b[25087] == 25087 && 
b[25088] == 25088 && 
b[25089] == 25089 && 
b[25090] == 25090 && 
b[25091] == 25091 && 
b[25092] == 25092 && 
b[25093] == 25093 && 
b[25094] == 25094 && 
b[25095] == 25095 && 
b[25096] == 25096 && 
b[25097] == 25097 && 
b[25098] == 25098 && 
b[25099] == 25099 && 
b[25100] == 25100 && 
b[25101] == 25101 && 
b[25102] == 25102 && 
b[25103] == 25103 && 
b[25104] == 25104 && 
b[25105] == 25105 && 
b[25106] == 25106 && 
b[25107] == 25107 && 
b[25108] == 25108 && 
b[25109] == 25109 && 
b[25110] == 25110 && 
b[25111] == 25111 && 
b[25112] == 25112 && 
b[25113] == 25113 && 
b[25114] == 25114 && 
b[25115] == 25115 && 
b[25116] == 25116 && 
b[25117] == 25117 && 
b[25118] == 25118 && 
b[25119] == 25119 && 
b[25120] == 25120 && 
b[25121] == 25121 && 
b[25122] == 25122 && 
b[25123] == 25123 && 
b[25124] == 25124 && 
b[25125] == 25125 && 
b[25126] == 25126 && 
b[25127] == 25127 && 
b[25128] == 25128 && 
b[25129] == 25129 && 
b[25130] == 25130 && 
b[25131] == 25131 && 
b[25132] == 25132 && 
b[25133] == 25133 && 
b[25134] == 25134 && 
b[25135] == 25135 && 
b[25136] == 25136 && 
b[25137] == 25137 && 
b[25138] == 25138 && 
b[25139] == 25139 && 
b[25140] == 25140 && 
b[25141] == 25141 && 
b[25142] == 25142 && 
b[25143] == 25143 && 
b[25144] == 25144 && 
b[25145] == 25145 && 
b[25146] == 25146 && 
b[25147] == 25147 && 
b[25148] == 25148 && 
b[25149] == 25149 && 
b[25150] == 25150 && 
b[25151] == 25151 && 
b[25152] == 25152 && 
b[25153] == 25153 && 
b[25154] == 25154 && 
b[25155] == 25155 && 
b[25156] == 25156 && 
b[25157] == 25157 && 
b[25158] == 25158 && 
b[25159] == 25159 && 
b[25160] == 25160 && 
b[25161] == 25161 && 
b[25162] == 25162 && 
b[25163] == 25163 && 
b[25164] == 25164 && 
b[25165] == 25165 && 
b[25166] == 25166 && 
b[25167] == 25167 && 
b[25168] == 25168 && 
b[25169] == 25169 && 
b[25170] == 25170 && 
b[25171] == 25171 && 
b[25172] == 25172 && 
b[25173] == 25173 && 
b[25174] == 25174 && 
b[25175] == 25175 && 
b[25176] == 25176 && 
b[25177] == 25177 && 
b[25178] == 25178 && 
b[25179] == 25179 && 
b[25180] == 25180 && 
b[25181] == 25181 && 
b[25182] == 25182 && 
b[25183] == 25183 && 
b[25184] == 25184 && 
b[25185] == 25185 && 
b[25186] == 25186 && 
b[25187] == 25187 && 
b[25188] == 25188 && 
b[25189] == 25189 && 
b[25190] == 25190 && 
b[25191] == 25191 && 
b[25192] == 25192 && 
b[25193] == 25193 && 
b[25194] == 25194 && 
b[25195] == 25195 && 
b[25196] == 25196 && 
b[25197] == 25197 && 
b[25198] == 25198 && 
b[25199] == 25199 && 
b[25200] == 25200 && 
b[25201] == 25201 && 
b[25202] == 25202 && 
b[25203] == 25203 && 
b[25204] == 25204 && 
b[25205] == 25205 && 
b[25206] == 25206 && 
b[25207] == 25207 && 
b[25208] == 25208 && 
b[25209] == 25209 && 
b[25210] == 25210 && 
b[25211] == 25211 && 
b[25212] == 25212 && 
b[25213] == 25213 && 
b[25214] == 25214 && 
b[25215] == 25215 && 
b[25216] == 25216 && 
b[25217] == 25217 && 
b[25218] == 25218 && 
b[25219] == 25219 && 
b[25220] == 25220 && 
b[25221] == 25221 && 
b[25222] == 25222 && 
b[25223] == 25223 && 
b[25224] == 25224 && 
b[25225] == 25225 && 
b[25226] == 25226 && 
b[25227] == 25227 && 
b[25228] == 25228 && 
b[25229] == 25229 && 
b[25230] == 25230 && 
b[25231] == 25231 && 
b[25232] == 25232 && 
b[25233] == 25233 && 
b[25234] == 25234 && 
b[25235] == 25235 && 
b[25236] == 25236 && 
b[25237] == 25237 && 
b[25238] == 25238 && 
b[25239] == 25239 && 
b[25240] == 25240 && 
b[25241] == 25241 && 
b[25242] == 25242 && 
b[25243] == 25243 && 
b[25244] == 25244 && 
b[25245] == 25245 && 
b[25246] == 25246 && 
b[25247] == 25247 && 
b[25248] == 25248 && 
b[25249] == 25249 && 
b[25250] == 25250 && 
b[25251] == 25251 && 
b[25252] == 25252 && 
b[25253] == 25253 && 
b[25254] == 25254 && 
b[25255] == 25255 && 
b[25256] == 25256 && 
b[25257] == 25257 && 
b[25258] == 25258 && 
b[25259] == 25259 && 
b[25260] == 25260 && 
b[25261] == 25261 && 
b[25262] == 25262 && 
b[25263] == 25263 && 
b[25264] == 25264 && 
b[25265] == 25265 && 
b[25266] == 25266 && 
b[25267] == 25267 && 
b[25268] == 25268 && 
b[25269] == 25269 && 
b[25270] == 25270 && 
b[25271] == 25271 && 
b[25272] == 25272 && 
b[25273] == 25273 && 
b[25274] == 25274 && 
b[25275] == 25275 && 
b[25276] == 25276 && 
b[25277] == 25277 && 
b[25278] == 25278 && 
b[25279] == 25279 && 
b[25280] == 25280 && 
b[25281] == 25281 && 
b[25282] == 25282 && 
b[25283] == 25283 && 
b[25284] == 25284 && 
b[25285] == 25285 && 
b[25286] == 25286 && 
b[25287] == 25287 && 
b[25288] == 25288 && 
b[25289] == 25289 && 
b[25290] == 25290 && 
b[25291] == 25291 && 
b[25292] == 25292 && 
b[25293] == 25293 && 
b[25294] == 25294 && 
b[25295] == 25295 && 
b[25296] == 25296 && 
b[25297] == 25297 && 
b[25298] == 25298 && 
b[25299] == 25299 && 
b[25300] == 25300 && 
b[25301] == 25301 && 
b[25302] == 25302 && 
b[25303] == 25303 && 
b[25304] == 25304 && 
b[25305] == 25305 && 
b[25306] == 25306 && 
b[25307] == 25307 && 
b[25308] == 25308 && 
b[25309] == 25309 && 
b[25310] == 25310 && 
b[25311] == 25311 && 
b[25312] == 25312 && 
b[25313] == 25313 && 
b[25314] == 25314 && 
b[25315] == 25315 && 
b[25316] == 25316 && 
b[25317] == 25317 && 
b[25318] == 25318 && 
b[25319] == 25319 && 
b[25320] == 25320 && 
b[25321] == 25321 && 
b[25322] == 25322 && 
b[25323] == 25323 && 
b[25324] == 25324 && 
b[25325] == 25325 && 
b[25326] == 25326 && 
b[25327] == 25327 && 
b[25328] == 25328 && 
b[25329] == 25329 && 
b[25330] == 25330 && 
b[25331] == 25331 && 
b[25332] == 25332 && 
b[25333] == 25333 && 
b[25334] == 25334 && 
b[25335] == 25335 && 
b[25336] == 25336 && 
b[25337] == 25337 && 
b[25338] == 25338 && 
b[25339] == 25339 && 
b[25340] == 25340 && 
b[25341] == 25341 && 
b[25342] == 25342 && 
b[25343] == 25343 && 
b[25344] == 25344 && 
b[25345] == 25345 && 
b[25346] == 25346 && 
b[25347] == 25347 && 
b[25348] == 25348 && 
b[25349] == 25349 && 
b[25350] == 25350 && 
b[25351] == 25351 && 
b[25352] == 25352 && 
b[25353] == 25353 && 
b[25354] == 25354 && 
b[25355] == 25355 && 
b[25356] == 25356 && 
b[25357] == 25357 && 
b[25358] == 25358 && 
b[25359] == 25359 && 
b[25360] == 25360 && 
b[25361] == 25361 && 
b[25362] == 25362 && 
b[25363] == 25363 && 
b[25364] == 25364 && 
b[25365] == 25365 && 
b[25366] == 25366 && 
b[25367] == 25367 && 
b[25368] == 25368 && 
b[25369] == 25369 && 
b[25370] == 25370 && 
b[25371] == 25371 && 
b[25372] == 25372 && 
b[25373] == 25373 && 
b[25374] == 25374 && 
b[25375] == 25375 && 
b[25376] == 25376 && 
b[25377] == 25377 && 
b[25378] == 25378 && 
b[25379] == 25379 && 
b[25380] == 25380 && 
b[25381] == 25381 && 
b[25382] == 25382 && 
b[25383] == 25383 && 
b[25384] == 25384 && 
b[25385] == 25385 && 
b[25386] == 25386 && 
b[25387] == 25387 && 
b[25388] == 25388 && 
b[25389] == 25389 && 
b[25390] == 25390 && 
b[25391] == 25391 && 
b[25392] == 25392 && 
b[25393] == 25393 && 
b[25394] == 25394 && 
b[25395] == 25395 && 
b[25396] == 25396 && 
b[25397] == 25397 && 
b[25398] == 25398 && 
b[25399] == 25399 && 
b[25400] == 25400 && 
b[25401] == 25401 && 
b[25402] == 25402 && 
b[25403] == 25403 && 
b[25404] == 25404 && 
b[25405] == 25405 && 
b[25406] == 25406 && 
b[25407] == 25407 && 
b[25408] == 25408 && 
b[25409] == 25409 && 
b[25410] == 25410 && 
b[25411] == 25411 && 
b[25412] == 25412 && 
b[25413] == 25413 && 
b[25414] == 25414 && 
b[25415] == 25415 && 
b[25416] == 25416 && 
b[25417] == 25417 && 
b[25418] == 25418 && 
b[25419] == 25419 && 
b[25420] == 25420 && 
b[25421] == 25421 && 
b[25422] == 25422 && 
b[25423] == 25423 && 
b[25424] == 25424 && 
b[25425] == 25425 && 
b[25426] == 25426 && 
b[25427] == 25427 && 
b[25428] == 25428 && 
b[25429] == 25429 && 
b[25430] == 25430 && 
b[25431] == 25431 && 
b[25432] == 25432 && 
b[25433] == 25433 && 
b[25434] == 25434 && 
b[25435] == 25435 && 
b[25436] == 25436 && 
b[25437] == 25437 && 
b[25438] == 25438 && 
b[25439] == 25439 && 
b[25440] == 25440 && 
b[25441] == 25441 && 
b[25442] == 25442 && 
b[25443] == 25443 && 
b[25444] == 25444 && 
b[25445] == 25445 && 
b[25446] == 25446 && 
b[25447] == 25447 && 
b[25448] == 25448 && 
b[25449] == 25449 && 
b[25450] == 25450 && 
b[25451] == 25451 && 
b[25452] == 25452 && 
b[25453] == 25453 && 
b[25454] == 25454 && 
b[25455] == 25455 && 
b[25456] == 25456 && 
b[25457] == 25457 && 
b[25458] == 25458 && 
b[25459] == 25459 && 
b[25460] == 25460 && 
b[25461] == 25461 && 
b[25462] == 25462 && 
b[25463] == 25463 && 
b[25464] == 25464 && 
b[25465] == 25465 && 
b[25466] == 25466 && 
b[25467] == 25467 && 
b[25468] == 25468 && 
b[25469] == 25469 && 
b[25470] == 25470 && 
b[25471] == 25471 && 
b[25472] == 25472 && 
b[25473] == 25473 && 
b[25474] == 25474 && 
b[25475] == 25475 && 
b[25476] == 25476 && 
b[25477] == 25477 && 
b[25478] == 25478 && 
b[25479] == 25479 && 
b[25480] == 25480 && 
b[25481] == 25481 && 
b[25482] == 25482 && 
b[25483] == 25483 && 
b[25484] == 25484 && 
b[25485] == 25485 && 
b[25486] == 25486 && 
b[25487] == 25487 && 
b[25488] == 25488 && 
b[25489] == 25489 && 
b[25490] == 25490 && 
b[25491] == 25491 && 
b[25492] == 25492 && 
b[25493] == 25493 && 
b[25494] == 25494 && 
b[25495] == 25495 && 
b[25496] == 25496 && 
b[25497] == 25497 && 
b[25498] == 25498 && 
b[25499] == 25499 && 
b[25500] == 25500 && 
b[25501] == 25501 && 
b[25502] == 25502 && 
b[25503] == 25503 && 
b[25504] == 25504 && 
b[25505] == 25505 && 
b[25506] == 25506 && 
b[25507] == 25507 && 
b[25508] == 25508 && 
b[25509] == 25509 && 
b[25510] == 25510 && 
b[25511] == 25511 && 
b[25512] == 25512 && 
b[25513] == 25513 && 
b[25514] == 25514 && 
b[25515] == 25515 && 
b[25516] == 25516 && 
b[25517] == 25517 && 
b[25518] == 25518 && 
b[25519] == 25519 && 
b[25520] == 25520 && 
b[25521] == 25521 && 
b[25522] == 25522 && 
b[25523] == 25523 && 
b[25524] == 25524 && 
b[25525] == 25525 && 
b[25526] == 25526 && 
b[25527] == 25527 && 
b[25528] == 25528 && 
b[25529] == 25529 && 
b[25530] == 25530 && 
b[25531] == 25531 && 
b[25532] == 25532 && 
b[25533] == 25533 && 
b[25534] == 25534 && 
b[25535] == 25535 && 
b[25536] == 25536 && 
b[25537] == 25537 && 
b[25538] == 25538 && 
b[25539] == 25539 && 
b[25540] == 25540 && 
b[25541] == 25541 && 
b[25542] == 25542 && 
b[25543] == 25543 && 
b[25544] == 25544 && 
b[25545] == 25545 && 
b[25546] == 25546 && 
b[25547] == 25547 && 
b[25548] == 25548 && 
b[25549] == 25549 && 
b[25550] == 25550 && 
b[25551] == 25551 && 
b[25552] == 25552 && 
b[25553] == 25553 && 
b[25554] == 25554 && 
b[25555] == 25555 && 
b[25556] == 25556 && 
b[25557] == 25557 && 
b[25558] == 25558 && 
b[25559] == 25559 && 
b[25560] == 25560 && 
b[25561] == 25561 && 
b[25562] == 25562 && 
b[25563] == 25563 && 
b[25564] == 25564 && 
b[25565] == 25565 && 
b[25566] == 25566 && 
b[25567] == 25567 && 
b[25568] == 25568 && 
b[25569] == 25569 && 
b[25570] == 25570 && 
b[25571] == 25571 && 
b[25572] == 25572 && 
b[25573] == 25573 && 
b[25574] == 25574 && 
b[25575] == 25575 && 
b[25576] == 25576 && 
b[25577] == 25577 && 
b[25578] == 25578 && 
b[25579] == 25579 && 
b[25580] == 25580 && 
b[25581] == 25581 && 
b[25582] == 25582 && 
b[25583] == 25583 && 
b[25584] == 25584 && 
b[25585] == 25585 && 
b[25586] == 25586 && 
b[25587] == 25587 && 
b[25588] == 25588 && 
b[25589] == 25589 && 
b[25590] == 25590 && 
b[25591] == 25591 && 
b[25592] == 25592 && 
b[25593] == 25593 && 
b[25594] == 25594 && 
b[25595] == 25595 && 
b[25596] == 25596 && 
b[25597] == 25597 && 
b[25598] == 25598 && 
b[25599] == 25599 && 
b[25600] == 25600 && 
b[25601] == 25601 && 
b[25602] == 25602 && 
b[25603] == 25603 && 
b[25604] == 25604 && 
b[25605] == 25605 && 
b[25606] == 25606 && 
b[25607] == 25607 && 
b[25608] == 25608 && 
b[25609] == 25609 && 
b[25610] == 25610 && 
b[25611] == 25611 && 
b[25612] == 25612 && 
b[25613] == 25613 && 
b[25614] == 25614 && 
b[25615] == 25615 && 
b[25616] == 25616 && 
b[25617] == 25617 && 
b[25618] == 25618 && 
b[25619] == 25619 && 
b[25620] == 25620 && 
b[25621] == 25621 && 
b[25622] == 25622 && 
b[25623] == 25623 && 
b[25624] == 25624 && 
b[25625] == 25625 && 
b[25626] == 25626 && 
b[25627] == 25627 && 
b[25628] == 25628 && 
b[25629] == 25629 && 
b[25630] == 25630 && 
b[25631] == 25631 && 
b[25632] == 25632 && 
b[25633] == 25633 && 
b[25634] == 25634 && 
b[25635] == 25635 && 
b[25636] == 25636 && 
b[25637] == 25637 && 
b[25638] == 25638 && 
b[25639] == 25639 && 
b[25640] == 25640 && 
b[25641] == 25641 && 
b[25642] == 25642 && 
b[25643] == 25643 && 
b[25644] == 25644 && 
b[25645] == 25645 && 
b[25646] == 25646 && 
b[25647] == 25647 && 
b[25648] == 25648 && 
b[25649] == 25649 && 
b[25650] == 25650 && 
b[25651] == 25651 && 
b[25652] == 25652 && 
b[25653] == 25653 && 
b[25654] == 25654 && 
b[25655] == 25655 && 
b[25656] == 25656 && 
b[25657] == 25657 && 
b[25658] == 25658 && 
b[25659] == 25659 && 
b[25660] == 25660 && 
b[25661] == 25661 && 
b[25662] == 25662 && 
b[25663] == 25663 && 
b[25664] == 25664 && 
b[25665] == 25665 && 
b[25666] == 25666 && 
b[25667] == 25667 && 
b[25668] == 25668 && 
b[25669] == 25669 && 
b[25670] == 25670 && 
b[25671] == 25671 && 
b[25672] == 25672 && 
b[25673] == 25673 && 
b[25674] == 25674 && 
b[25675] == 25675 && 
b[25676] == 25676 && 
b[25677] == 25677 && 
b[25678] == 25678 && 
b[25679] == 25679 && 
b[25680] == 25680 && 
b[25681] == 25681 && 
b[25682] == 25682 && 
b[25683] == 25683 && 
b[25684] == 25684 && 
b[25685] == 25685 && 
b[25686] == 25686 && 
b[25687] == 25687 && 
b[25688] == 25688 && 
b[25689] == 25689 && 
b[25690] == 25690 && 
b[25691] == 25691 && 
b[25692] == 25692 && 
b[25693] == 25693 && 
b[25694] == 25694 && 
b[25695] == 25695 && 
b[25696] == 25696 && 
b[25697] == 25697 && 
b[25698] == 25698 && 
b[25699] == 25699 && 
b[25700] == 25700 && 
b[25701] == 25701 && 
b[25702] == 25702 && 
b[25703] == 25703 && 
b[25704] == 25704 && 
b[25705] == 25705 && 
b[25706] == 25706 && 
b[25707] == 25707 && 
b[25708] == 25708 && 
b[25709] == 25709 && 
b[25710] == 25710 && 
b[25711] == 25711 && 
b[25712] == 25712 && 
b[25713] == 25713 && 
b[25714] == 25714 && 
b[25715] == 25715 && 
b[25716] == 25716 && 
b[25717] == 25717 && 
b[25718] == 25718 && 
b[25719] == 25719 && 
b[25720] == 25720 && 
b[25721] == 25721 && 
b[25722] == 25722 && 
b[25723] == 25723 && 
b[25724] == 25724 && 
b[25725] == 25725 && 
b[25726] == 25726 && 
b[25727] == 25727 && 
b[25728] == 25728 && 
b[25729] == 25729 && 
b[25730] == 25730 && 
b[25731] == 25731 && 
b[25732] == 25732 && 
b[25733] == 25733 && 
b[25734] == 25734 && 
b[25735] == 25735 && 
b[25736] == 25736 && 
b[25737] == 25737 && 
b[25738] == 25738 && 
b[25739] == 25739 && 
b[25740] == 25740 && 
b[25741] == 25741 && 
b[25742] == 25742 && 
b[25743] == 25743 && 
b[25744] == 25744 && 
b[25745] == 25745 && 
b[25746] == 25746 && 
b[25747] == 25747 && 
b[25748] == 25748 && 
b[25749] == 25749 && 
b[25750] == 25750 && 
b[25751] == 25751 && 
b[25752] == 25752 && 
b[25753] == 25753 && 
b[25754] == 25754 && 
b[25755] == 25755 && 
b[25756] == 25756 && 
b[25757] == 25757 && 
b[25758] == 25758 && 
b[25759] == 25759 && 
b[25760] == 25760 && 
b[25761] == 25761 && 
b[25762] == 25762 && 
b[25763] == 25763 && 
b[25764] == 25764 && 
b[25765] == 25765 && 
b[25766] == 25766 && 
b[25767] == 25767 && 
b[25768] == 25768 && 
b[25769] == 25769 && 
b[25770] == 25770 && 
b[25771] == 25771 && 
b[25772] == 25772 && 
b[25773] == 25773 && 
b[25774] == 25774 && 
b[25775] == 25775 && 
b[25776] == 25776 && 
b[25777] == 25777 && 
b[25778] == 25778 && 
b[25779] == 25779 && 
b[25780] == 25780 && 
b[25781] == 25781 && 
b[25782] == 25782 && 
b[25783] == 25783 && 
b[25784] == 25784 && 
b[25785] == 25785 && 
b[25786] == 25786 && 
b[25787] == 25787 && 
b[25788] == 25788 && 
b[25789] == 25789 && 
b[25790] == 25790 && 
b[25791] == 25791 && 
b[25792] == 25792 && 
b[25793] == 25793 && 
b[25794] == 25794 && 
b[25795] == 25795 && 
b[25796] == 25796 && 
b[25797] == 25797 && 
b[25798] == 25798 && 
b[25799] == 25799 && 
b[25800] == 25800 && 
b[25801] == 25801 && 
b[25802] == 25802 && 
b[25803] == 25803 && 
b[25804] == 25804 && 
b[25805] == 25805 && 
b[25806] == 25806 && 
b[25807] == 25807 && 
b[25808] == 25808 && 
b[25809] == 25809 && 
b[25810] == 25810 && 
b[25811] == 25811 && 
b[25812] == 25812 && 
b[25813] == 25813 && 
b[25814] == 25814 && 
b[25815] == 25815 && 
b[25816] == 25816 && 
b[25817] == 25817 && 
b[25818] == 25818 && 
b[25819] == 25819 && 
b[25820] == 25820 && 
b[25821] == 25821 && 
b[25822] == 25822 && 
b[25823] == 25823 && 
b[25824] == 25824 && 
b[25825] == 25825 && 
b[25826] == 25826 && 
b[25827] == 25827 && 
b[25828] == 25828 && 
b[25829] == 25829 && 
b[25830] == 25830 && 
b[25831] == 25831 && 
b[25832] == 25832 && 
b[25833] == 25833 && 
b[25834] == 25834 && 
b[25835] == 25835 && 
b[25836] == 25836 && 
b[25837] == 25837 && 
b[25838] == 25838 && 
b[25839] == 25839 && 
b[25840] == 25840 && 
b[25841] == 25841 && 
b[25842] == 25842 && 
b[25843] == 25843 && 
b[25844] == 25844 && 
b[25845] == 25845 && 
b[25846] == 25846 && 
b[25847] == 25847 && 
b[25848] == 25848 && 
b[25849] == 25849 && 
b[25850] == 25850 && 
b[25851] == 25851 && 
b[25852] == 25852 && 
b[25853] == 25853 && 
b[25854] == 25854 && 
b[25855] == 25855 && 
b[25856] == 25856 && 
b[25857] == 25857 && 
b[25858] == 25858 && 
b[25859] == 25859 && 
b[25860] == 25860 && 
b[25861] == 25861 && 
b[25862] == 25862 && 
b[25863] == 25863 && 
b[25864] == 25864 && 
b[25865] == 25865 && 
b[25866] == 25866 && 
b[25867] == 25867 && 
b[25868] == 25868 && 
b[25869] == 25869 && 
b[25870] == 25870 && 
b[25871] == 25871 && 
b[25872] == 25872 && 
b[25873] == 25873 && 
b[25874] == 25874 && 
b[25875] == 25875 && 
b[25876] == 25876 && 
b[25877] == 25877 && 
b[25878] == 25878 && 
b[25879] == 25879 && 
b[25880] == 25880 && 
b[25881] == 25881 && 
b[25882] == 25882 && 
b[25883] == 25883 && 
b[25884] == 25884 && 
b[25885] == 25885 && 
b[25886] == 25886 && 
b[25887] == 25887 && 
b[25888] == 25888 && 
b[25889] == 25889 && 
b[25890] == 25890 && 
b[25891] == 25891 && 
b[25892] == 25892 && 
b[25893] == 25893 && 
b[25894] == 25894 && 
b[25895] == 25895 && 
b[25896] == 25896 && 
b[25897] == 25897 && 
b[25898] == 25898 && 
b[25899] == 25899 && 
b[25900] == 25900 && 
b[25901] == 25901 && 
b[25902] == 25902 && 
b[25903] == 25903 && 
b[25904] == 25904 && 
b[25905] == 25905 && 
b[25906] == 25906 && 
b[25907] == 25907 && 
b[25908] == 25908 && 
b[25909] == 25909 && 
b[25910] == 25910 && 
b[25911] == 25911 && 
b[25912] == 25912 && 
b[25913] == 25913 && 
b[25914] == 25914 && 
b[25915] == 25915 && 
b[25916] == 25916 && 
b[25917] == 25917 && 
b[25918] == 25918 && 
b[25919] == 25919 && 
b[25920] == 25920 && 
b[25921] == 25921 && 
b[25922] == 25922 && 
b[25923] == 25923 && 
b[25924] == 25924 && 
b[25925] == 25925 && 
b[25926] == 25926 && 
b[25927] == 25927 && 
b[25928] == 25928 && 
b[25929] == 25929 && 
b[25930] == 25930 && 
b[25931] == 25931 && 
b[25932] == 25932 && 
b[25933] == 25933 && 
b[25934] == 25934 && 
b[25935] == 25935 && 
b[25936] == 25936 && 
b[25937] == 25937 && 
b[25938] == 25938 && 
b[25939] == 25939 && 
b[25940] == 25940 && 
b[25941] == 25941 && 
b[25942] == 25942 && 
b[25943] == 25943 && 
b[25944] == 25944 && 
b[25945] == 25945 && 
b[25946] == 25946 && 
b[25947] == 25947 && 
b[25948] == 25948 && 
b[25949] == 25949 && 
b[25950] == 25950 && 
b[25951] == 25951 && 
b[25952] == 25952 && 
b[25953] == 25953 && 
b[25954] == 25954 && 
b[25955] == 25955 && 
b[25956] == 25956 && 
b[25957] == 25957 && 
b[25958] == 25958 && 
b[25959] == 25959 && 
b[25960] == 25960 && 
b[25961] == 25961 && 
b[25962] == 25962 && 
b[25963] == 25963 && 
b[25964] == 25964 && 
b[25965] == 25965 && 
b[25966] == 25966 && 
b[25967] == 25967 && 
b[25968] == 25968 && 
b[25969] == 25969 && 
b[25970] == 25970 && 
b[25971] == 25971 && 
b[25972] == 25972 && 
b[25973] == 25973 && 
b[25974] == 25974 && 
b[25975] == 25975 && 
b[25976] == 25976 && 
b[25977] == 25977 && 
b[25978] == 25978 && 
b[25979] == 25979 && 
b[25980] == 25980 && 
b[25981] == 25981 && 
b[25982] == 25982 && 
b[25983] == 25983 && 
b[25984] == 25984 && 
b[25985] == 25985 && 
b[25986] == 25986 && 
b[25987] == 25987 && 
b[25988] == 25988 && 
b[25989] == 25989 && 
b[25990] == 25990 && 
b[25991] == 25991 && 
b[25992] == 25992 && 
b[25993] == 25993 && 
b[25994] == 25994 && 
b[25995] == 25995 && 
b[25996] == 25996 && 
b[25997] == 25997 && 
b[25998] == 25998 && 
b[25999] == 25999 && 
b[26000] == 26000 && 
b[26001] == 26001 && 
b[26002] == 26002 && 
b[26003] == 26003 && 
b[26004] == 26004 && 
b[26005] == 26005 && 
b[26006] == 26006 && 
b[26007] == 26007 && 
b[26008] == 26008 && 
b[26009] == 26009 && 
b[26010] == 26010 && 
b[26011] == 26011 && 
b[26012] == 26012 && 
b[26013] == 26013 && 
b[26014] == 26014 && 
b[26015] == 26015 && 
b[26016] == 26016 && 
b[26017] == 26017 && 
b[26018] == 26018 && 
b[26019] == 26019 && 
b[26020] == 26020 && 
b[26021] == 26021 && 
b[26022] == 26022 && 
b[26023] == 26023 && 
b[26024] == 26024 && 
b[26025] == 26025 && 
b[26026] == 26026 && 
b[26027] == 26027 && 
b[26028] == 26028 && 
b[26029] == 26029 && 
b[26030] == 26030 && 
b[26031] == 26031 && 
b[26032] == 26032 && 
b[26033] == 26033 && 
b[26034] == 26034 && 
b[26035] == 26035 && 
b[26036] == 26036 && 
b[26037] == 26037 && 
b[26038] == 26038 && 
b[26039] == 26039 && 
b[26040] == 26040 && 
b[26041] == 26041 && 
b[26042] == 26042 && 
b[26043] == 26043 && 
b[26044] == 26044 && 
b[26045] == 26045 && 
b[26046] == 26046 && 
b[26047] == 26047 && 
b[26048] == 26048 && 
b[26049] == 26049 && 
b[26050] == 26050 && 
b[26051] == 26051 && 
b[26052] == 26052 && 
b[26053] == 26053 && 
b[26054] == 26054 && 
b[26055] == 26055 && 
b[26056] == 26056 && 
b[26057] == 26057 && 
b[26058] == 26058 && 
b[26059] == 26059 && 
b[26060] == 26060 && 
b[26061] == 26061 && 
b[26062] == 26062 && 
b[26063] == 26063 && 
b[26064] == 26064 && 
b[26065] == 26065 && 
b[26066] == 26066 && 
b[26067] == 26067 && 
b[26068] == 26068 && 
b[26069] == 26069 && 
b[26070] == 26070 && 
b[26071] == 26071 && 
b[26072] == 26072 && 
b[26073] == 26073 && 
b[26074] == 26074 && 
b[26075] == 26075 && 
b[26076] == 26076 && 
b[26077] == 26077 && 
b[26078] == 26078 && 
b[26079] == 26079 && 
b[26080] == 26080 && 
b[26081] == 26081 && 
b[26082] == 26082 && 
b[26083] == 26083 && 
b[26084] == 26084 && 
b[26085] == 26085 && 
b[26086] == 26086 && 
b[26087] == 26087 && 
b[26088] == 26088 && 
b[26089] == 26089 && 
b[26090] == 26090 && 
b[26091] == 26091 && 
b[26092] == 26092 && 
b[26093] == 26093 && 
b[26094] == 26094 && 
b[26095] == 26095 && 
b[26096] == 26096 && 
b[26097] == 26097 && 
b[26098] == 26098 && 
b[26099] == 26099 && 
b[26100] == 26100 && 
b[26101] == 26101 && 
b[26102] == 26102 && 
b[26103] == 26103 && 
b[26104] == 26104 && 
b[26105] == 26105 && 
b[26106] == 26106 && 
b[26107] == 26107 && 
b[26108] == 26108 && 
b[26109] == 26109 && 
b[26110] == 26110 && 
b[26111] == 26111 && 
b[26112] == 26112 && 
b[26113] == 26113 && 
b[26114] == 26114 && 
b[26115] == 26115 && 
b[26116] == 26116 && 
b[26117] == 26117 && 
b[26118] == 26118 && 
b[26119] == 26119 && 
b[26120] == 26120 && 
b[26121] == 26121 && 
b[26122] == 26122 && 
b[26123] == 26123 && 
b[26124] == 26124 && 
b[26125] == 26125 && 
b[26126] == 26126 && 
b[26127] == 26127 && 
b[26128] == 26128 && 
b[26129] == 26129 && 
b[26130] == 26130 && 
b[26131] == 26131 && 
b[26132] == 26132 && 
b[26133] == 26133 && 
b[26134] == 26134 && 
b[26135] == 26135 && 
b[26136] == 26136 && 
b[26137] == 26137 && 
b[26138] == 26138 && 
b[26139] == 26139 && 
b[26140] == 26140 && 
b[26141] == 26141 && 
b[26142] == 26142 && 
b[26143] == 26143 && 
b[26144] == 26144 && 
b[26145] == 26145 && 
b[26146] == 26146 && 
b[26147] == 26147 && 
b[26148] == 26148 && 
b[26149] == 26149 && 
b[26150] == 26150 && 
b[26151] == 26151 && 
b[26152] == 26152 && 
b[26153] == 26153 && 
b[26154] == 26154 && 
b[26155] == 26155 && 
b[26156] == 26156 && 
b[26157] == 26157 && 
b[26158] == 26158 && 
b[26159] == 26159 && 
b[26160] == 26160 && 
b[26161] == 26161 && 
b[26162] == 26162 && 
b[26163] == 26163 && 
b[26164] == 26164 && 
b[26165] == 26165 && 
b[26166] == 26166 && 
b[26167] == 26167 && 
b[26168] == 26168 && 
b[26169] == 26169 && 
b[26170] == 26170 && 
b[26171] == 26171 && 
b[26172] == 26172 && 
b[26173] == 26173 && 
b[26174] == 26174 && 
b[26175] == 26175 && 
b[26176] == 26176 && 
b[26177] == 26177 && 
b[26178] == 26178 && 
b[26179] == 26179 && 
b[26180] == 26180 && 
b[26181] == 26181 && 
b[26182] == 26182 && 
b[26183] == 26183 && 
b[26184] == 26184 && 
b[26185] == 26185 && 
b[26186] == 26186 && 
b[26187] == 26187 && 
b[26188] == 26188 && 
b[26189] == 26189 && 
b[26190] == 26190 && 
b[26191] == 26191 && 
b[26192] == 26192 && 
b[26193] == 26193 && 
b[26194] == 26194 && 
b[26195] == 26195 && 
b[26196] == 26196 && 
b[26197] == 26197 && 
b[26198] == 26198 && 
b[26199] == 26199 && 
b[26200] == 26200 && 
b[26201] == 26201 && 
b[26202] == 26202 && 
b[26203] == 26203 && 
b[26204] == 26204 && 
b[26205] == 26205 && 
b[26206] == 26206 && 
b[26207] == 26207 && 
b[26208] == 26208 && 
b[26209] == 26209 && 
b[26210] == 26210 && 
b[26211] == 26211 && 
b[26212] == 26212 && 
b[26213] == 26213 && 
b[26214] == 26214 && 
b[26215] == 26215 && 
b[26216] == 26216 && 
b[26217] == 26217 && 
b[26218] == 26218 && 
b[26219] == 26219 && 
b[26220] == 26220 && 
b[26221] == 26221 && 
b[26222] == 26222 && 
b[26223] == 26223 && 
b[26224] == 26224 && 
b[26225] == 26225 && 
b[26226] == 26226 && 
b[26227] == 26227 && 
b[26228] == 26228 && 
b[26229] == 26229 && 
b[26230] == 26230 && 
b[26231] == 26231 && 
b[26232] == 26232 && 
b[26233] == 26233 && 
b[26234] == 26234 && 
b[26235] == 26235 && 
b[26236] == 26236 && 
b[26237] == 26237 && 
b[26238] == 26238 && 
b[26239] == 26239 && 
b[26240] == 26240 && 
b[26241] == 26241 && 
b[26242] == 26242 && 
b[26243] == 26243 && 
b[26244] == 26244 && 
b[26245] == 26245 && 
b[26246] == 26246 && 
b[26247] == 26247 && 
b[26248] == 26248 && 
b[26249] == 26249 && 
b[26250] == 26250 && 
b[26251] == 26251 && 
b[26252] == 26252 && 
b[26253] == 26253 && 
b[26254] == 26254 && 
b[26255] == 26255 && 
b[26256] == 26256 && 
b[26257] == 26257 && 
b[26258] == 26258 && 
b[26259] == 26259 && 
b[26260] == 26260 && 
b[26261] == 26261 && 
b[26262] == 26262 && 
b[26263] == 26263 && 
b[26264] == 26264 && 
b[26265] == 26265 && 
b[26266] == 26266 && 
b[26267] == 26267 && 
b[26268] == 26268 && 
b[26269] == 26269 && 
b[26270] == 26270 && 
b[26271] == 26271 && 
b[26272] == 26272 && 
b[26273] == 26273 && 
b[26274] == 26274 && 
b[26275] == 26275 && 
b[26276] == 26276 && 
b[26277] == 26277 && 
b[26278] == 26278 && 
b[26279] == 26279 && 
b[26280] == 26280 && 
b[26281] == 26281 && 
b[26282] == 26282 && 
b[26283] == 26283 && 
b[26284] == 26284 && 
b[26285] == 26285 && 
b[26286] == 26286 && 
b[26287] == 26287 && 
b[26288] == 26288 && 
b[26289] == 26289 && 
b[26290] == 26290 && 
b[26291] == 26291 && 
b[26292] == 26292 && 
b[26293] == 26293 && 
b[26294] == 26294 && 
b[26295] == 26295 && 
b[26296] == 26296 && 
b[26297] == 26297 && 
b[26298] == 26298 && 
b[26299] == 26299 && 
b[26300] == 26300 && 
b[26301] == 26301 && 
b[26302] == 26302 && 
b[26303] == 26303 && 
b[26304] == 26304 && 
b[26305] == 26305 && 
b[26306] == 26306 && 
b[26307] == 26307 && 
b[26308] == 26308 && 
b[26309] == 26309 && 
b[26310] == 26310 && 
b[26311] == 26311 && 
b[26312] == 26312 && 
b[26313] == 26313 && 
b[26314] == 26314 && 
b[26315] == 26315 && 
b[26316] == 26316 && 
b[26317] == 26317 && 
b[26318] == 26318 && 
b[26319] == 26319 && 
b[26320] == 26320 && 
b[26321] == 26321 && 
b[26322] == 26322 && 
b[26323] == 26323 && 
b[26324] == 26324 && 
b[26325] == 26325 && 
b[26326] == 26326 && 
b[26327] == 26327 && 
b[26328] == 26328 && 
b[26329] == 26329 && 
b[26330] == 26330 && 
b[26331] == 26331 && 
b[26332] == 26332 && 
b[26333] == 26333 && 
b[26334] == 26334 && 
b[26335] == 26335 && 
b[26336] == 26336 && 
b[26337] == 26337 && 
b[26338] == 26338 && 
b[26339] == 26339 && 
b[26340] == 26340 && 
b[26341] == 26341 && 
b[26342] == 26342 && 
b[26343] == 26343 && 
b[26344] == 26344 && 
b[26345] == 26345 && 
b[26346] == 26346 && 
b[26347] == 26347 && 
b[26348] == 26348 && 
b[26349] == 26349 && 
b[26350] == 26350 && 
b[26351] == 26351 && 
b[26352] == 26352 && 
b[26353] == 26353 && 
b[26354] == 26354 && 
b[26355] == 26355 && 
b[26356] == 26356 && 
b[26357] == 26357 && 
b[26358] == 26358 && 
b[26359] == 26359 && 
b[26360] == 26360 && 
b[26361] == 26361 && 
b[26362] == 26362 && 
b[26363] == 26363 && 
b[26364] == 26364 && 
b[26365] == 26365 && 
b[26366] == 26366 && 
b[26367] == 26367 && 
b[26368] == 26368 && 
b[26369] == 26369 && 
b[26370] == 26370 && 
b[26371] == 26371 && 
b[26372] == 26372 && 
b[26373] == 26373 && 
b[26374] == 26374 && 
b[26375] == 26375 && 
b[26376] == 26376 && 
b[26377] == 26377 && 
b[26378] == 26378 && 
b[26379] == 26379 && 
b[26380] == 26380 && 
b[26381] == 26381 && 
b[26382] == 26382 && 
b[26383] == 26383 && 
b[26384] == 26384 && 
b[26385] == 26385 && 
b[26386] == 26386 && 
b[26387] == 26387 && 
b[26388] == 26388 && 
b[26389] == 26389 && 
b[26390] == 26390 && 
b[26391] == 26391 && 
b[26392] == 26392 && 
b[26393] == 26393 && 
b[26394] == 26394 && 
b[26395] == 26395 && 
b[26396] == 26396 && 
b[26397] == 26397 && 
b[26398] == 26398 && 
b[26399] == 26399 && 
b[26400] == 26400 && 
b[26401] == 26401 && 
b[26402] == 26402 && 
b[26403] == 26403 && 
b[26404] == 26404 && 
b[26405] == 26405 && 
b[26406] == 26406 && 
b[26407] == 26407 && 
b[26408] == 26408 && 
b[26409] == 26409 && 
b[26410] == 26410 && 
b[26411] == 26411 && 
b[26412] == 26412 && 
b[26413] == 26413 && 
b[26414] == 26414 && 
b[26415] == 26415 && 
b[26416] == 26416 && 
b[26417] == 26417 && 
b[26418] == 26418 && 
b[26419] == 26419 && 
b[26420] == 26420 && 
b[26421] == 26421 && 
b[26422] == 26422 && 
b[26423] == 26423 && 
b[26424] == 26424 && 
b[26425] == 26425 && 
b[26426] == 26426 && 
b[26427] == 26427 && 
b[26428] == 26428 && 
b[26429] == 26429 && 
b[26430] == 26430 && 
b[26431] == 26431 && 
b[26432] == 26432 && 
b[26433] == 26433 && 
b[26434] == 26434 && 
b[26435] == 26435 && 
b[26436] == 26436 && 
b[26437] == 26437 && 
b[26438] == 26438 && 
b[26439] == 26439 && 
b[26440] == 26440 && 
b[26441] == 26441 && 
b[26442] == 26442 && 
b[26443] == 26443 && 
b[26444] == 26444 && 
b[26445] == 26445 && 
b[26446] == 26446 && 
b[26447] == 26447 && 
b[26448] == 26448 && 
b[26449] == 26449 && 
b[26450] == 26450 && 
b[26451] == 26451 && 
b[26452] == 26452 && 
b[26453] == 26453 && 
b[26454] == 26454 && 
b[26455] == 26455 && 
b[26456] == 26456 && 
b[26457] == 26457 && 
b[26458] == 26458 && 
b[26459] == 26459 && 
b[26460] == 26460 && 
b[26461] == 26461 && 
b[26462] == 26462 && 
b[26463] == 26463 && 
b[26464] == 26464 && 
b[26465] == 26465 && 
b[26466] == 26466 && 
b[26467] == 26467 && 
b[26468] == 26468 && 
b[26469] == 26469 && 
b[26470] == 26470 && 
b[26471] == 26471 && 
b[26472] == 26472 && 
b[26473] == 26473 && 
b[26474] == 26474 && 
b[26475] == 26475 && 
b[26476] == 26476 && 
b[26477] == 26477 && 
b[26478] == 26478 && 
b[26479] == 26479 && 
b[26480] == 26480 && 
b[26481] == 26481 && 
b[26482] == 26482 && 
b[26483] == 26483 && 
b[26484] == 26484 && 
b[26485] == 26485 && 
b[26486] == 26486 && 
b[26487] == 26487 && 
b[26488] == 26488 && 
b[26489] == 26489 && 
b[26490] == 26490 && 
b[26491] == 26491 && 
b[26492] == 26492 && 
b[26493] == 26493 && 
b[26494] == 26494 && 
b[26495] == 26495 && 
b[26496] == 26496 && 
b[26497] == 26497 && 
b[26498] == 26498 && 
b[26499] == 26499 && 
b[26500] == 26500 && 
b[26501] == 26501 && 
b[26502] == 26502 && 
b[26503] == 26503 && 
b[26504] == 26504 && 
b[26505] == 26505 && 
b[26506] == 26506 && 
b[26507] == 26507 && 
b[26508] == 26508 && 
b[26509] == 26509 && 
b[26510] == 26510 && 
b[26511] == 26511 && 
b[26512] == 26512 && 
b[26513] == 26513 && 
b[26514] == 26514 && 
b[26515] == 26515 && 
b[26516] == 26516 && 
b[26517] == 26517 && 
b[26518] == 26518 && 
b[26519] == 26519 && 
b[26520] == 26520 && 
b[26521] == 26521 && 
b[26522] == 26522 && 
b[26523] == 26523 && 
b[26524] == 26524 && 
b[26525] == 26525 && 
b[26526] == 26526 && 
b[26527] == 26527 && 
b[26528] == 26528 && 
b[26529] == 26529 && 
b[26530] == 26530 && 
b[26531] == 26531 && 
b[26532] == 26532 && 
b[26533] == 26533 && 
b[26534] == 26534 && 
b[26535] == 26535 && 
b[26536] == 26536 && 
b[26537] == 26537 && 
b[26538] == 26538 && 
b[26539] == 26539 && 
b[26540] == 26540 && 
b[26541] == 26541 && 
b[26542] == 26542 && 
b[26543] == 26543 && 
b[26544] == 26544 && 
b[26545] == 26545 && 
b[26546] == 26546 && 
b[26547] == 26547 && 
b[26548] == 26548 && 
b[26549] == 26549 && 
b[26550] == 26550 && 
b[26551] == 26551 && 
b[26552] == 26552 && 
b[26553] == 26553 && 
b[26554] == 26554 && 
b[26555] == 26555 && 
b[26556] == 26556 && 
b[26557] == 26557 && 
b[26558] == 26558 && 
b[26559] == 26559 && 
b[26560] == 26560 && 
b[26561] == 26561 && 
b[26562] == 26562 && 
b[26563] == 26563 && 
b[26564] == 26564 && 
b[26565] == 26565 && 
b[26566] == 26566 && 
b[26567] == 26567 && 
b[26568] == 26568 && 
b[26569] == 26569 && 
b[26570] == 26570 && 
b[26571] == 26571 && 
b[26572] == 26572 && 
b[26573] == 26573 && 
b[26574] == 26574 && 
b[26575] == 26575 && 
b[26576] == 26576 && 
b[26577] == 26577 && 
b[26578] == 26578 && 
b[26579] == 26579 && 
b[26580] == 26580 && 
b[26581] == 26581 && 
b[26582] == 26582 && 
b[26583] == 26583 && 
b[26584] == 26584 && 
b[26585] == 26585 && 
b[26586] == 26586 && 
b[26587] == 26587 && 
b[26588] == 26588 && 
b[26589] == 26589 && 
b[26590] == 26590 && 
b[26591] == 26591 && 
b[26592] == 26592 && 
b[26593] == 26593 && 
b[26594] == 26594 && 
b[26595] == 26595 && 
b[26596] == 26596 && 
b[26597] == 26597 && 
b[26598] == 26598 && 
b[26599] == 26599 && 
b[26600] == 26600 && 
b[26601] == 26601 && 
b[26602] == 26602 && 
b[26603] == 26603 && 
b[26604] == 26604 && 
b[26605] == 26605 && 
b[26606] == 26606 && 
b[26607] == 26607 && 
b[26608] == 26608 && 
b[26609] == 26609 && 
b[26610] == 26610 && 
b[26611] == 26611 && 
b[26612] == 26612 && 
b[26613] == 26613 && 
b[26614] == 26614 && 
b[26615] == 26615 && 
b[26616] == 26616 && 
b[26617] == 26617 && 
b[26618] == 26618 && 
b[26619] == 26619 && 
b[26620] == 26620 && 
b[26621] == 26621 && 
b[26622] == 26622 && 
b[26623] == 26623 && 
b[26624] == 26624 && 
b[26625] == 26625 && 
b[26626] == 26626 && 
b[26627] == 26627 && 
b[26628] == 26628 && 
b[26629] == 26629 && 
b[26630] == 26630 && 
b[26631] == 26631 && 
b[26632] == 26632 && 
b[26633] == 26633 && 
b[26634] == 26634 && 
b[26635] == 26635 && 
b[26636] == 26636 && 
b[26637] == 26637 && 
b[26638] == 26638 && 
b[26639] == 26639 && 
b[26640] == 26640 && 
b[26641] == 26641 && 
b[26642] == 26642 && 
b[26643] == 26643 && 
b[26644] == 26644 && 
b[26645] == 26645 && 
b[26646] == 26646 && 
b[26647] == 26647 && 
b[26648] == 26648 && 
b[26649] == 26649 && 
b[26650] == 26650 && 
b[26651] == 26651 && 
b[26652] == 26652 && 
b[26653] == 26653 && 
b[26654] == 26654 && 
b[26655] == 26655 && 
b[26656] == 26656 && 
b[26657] == 26657 && 
b[26658] == 26658 && 
b[26659] == 26659 && 
b[26660] == 26660 && 
b[26661] == 26661 && 
b[26662] == 26662 && 
b[26663] == 26663 && 
b[26664] == 26664 && 
b[26665] == 26665 && 
b[26666] == 26666 && 
b[26667] == 26667 && 
b[26668] == 26668 && 
b[26669] == 26669 && 
b[26670] == 26670 && 
b[26671] == 26671 && 
b[26672] == 26672 && 
b[26673] == 26673 && 
b[26674] == 26674 && 
b[26675] == 26675 && 
b[26676] == 26676 && 
b[26677] == 26677 && 
b[26678] == 26678 && 
b[26679] == 26679 && 
b[26680] == 26680 && 
b[26681] == 26681 && 
b[26682] == 26682 && 
b[26683] == 26683 && 
b[26684] == 26684 && 
b[26685] == 26685 && 
b[26686] == 26686 && 
b[26687] == 26687 && 
b[26688] == 26688 && 
b[26689] == 26689 && 
b[26690] == 26690 && 
b[26691] == 26691 && 
b[26692] == 26692 && 
b[26693] == 26693 && 
b[26694] == 26694 && 
b[26695] == 26695 && 
b[26696] == 26696 && 
b[26697] == 26697 && 
b[26698] == 26698 && 
b[26699] == 26699 && 
b[26700] == 26700 && 
b[26701] == 26701 && 
b[26702] == 26702 && 
b[26703] == 26703 && 
b[26704] == 26704 && 
b[26705] == 26705 && 
b[26706] == 26706 && 
b[26707] == 26707 && 
b[26708] == 26708 && 
b[26709] == 26709 && 
b[26710] == 26710 && 
b[26711] == 26711 && 
b[26712] == 26712 && 
b[26713] == 26713 && 
b[26714] == 26714 && 
b[26715] == 26715 && 
b[26716] == 26716 && 
b[26717] == 26717 && 
b[26718] == 26718 && 
b[26719] == 26719 && 
b[26720] == 26720 && 
b[26721] == 26721 && 
b[26722] == 26722 && 
b[26723] == 26723 && 
b[26724] == 26724 && 
b[26725] == 26725 && 
b[26726] == 26726 && 
b[26727] == 26727 && 
b[26728] == 26728 && 
b[26729] == 26729 && 
b[26730] == 26730 && 
b[26731] == 26731 && 
b[26732] == 26732 && 
b[26733] == 26733 && 
b[26734] == 26734 && 
b[26735] == 26735 && 
b[26736] == 26736 && 
b[26737] == 26737 && 
b[26738] == 26738 && 
b[26739] == 26739 && 
b[26740] == 26740 && 
b[26741] == 26741 && 
b[26742] == 26742 && 
b[26743] == 26743 && 
b[26744] == 26744 && 
b[26745] == 26745 && 
b[26746] == 26746 && 
b[26747] == 26747 && 
b[26748] == 26748 && 
b[26749] == 26749 && 
b[26750] == 26750 && 
b[26751] == 26751 && 
b[26752] == 26752 && 
b[26753] == 26753 && 
b[26754] == 26754 && 
b[26755] == 26755 && 
b[26756] == 26756 && 
b[26757] == 26757 && 
b[26758] == 26758 && 
b[26759] == 26759 && 
b[26760] == 26760 && 
b[26761] == 26761 && 
b[26762] == 26762 && 
b[26763] == 26763 && 
b[26764] == 26764 && 
b[26765] == 26765 && 
b[26766] == 26766 && 
b[26767] == 26767 && 
b[26768] == 26768 && 
b[26769] == 26769 && 
b[26770] == 26770 && 
b[26771] == 26771 && 
b[26772] == 26772 && 
b[26773] == 26773 && 
b[26774] == 26774 && 
b[26775] == 26775 && 
b[26776] == 26776 && 
b[26777] == 26777 && 
b[26778] == 26778 && 
b[26779] == 26779 && 
b[26780] == 26780 && 
b[26781] == 26781 && 
b[26782] == 26782 && 
b[26783] == 26783 && 
b[26784] == 26784 && 
b[26785] == 26785 && 
b[26786] == 26786 && 
b[26787] == 26787 && 
b[26788] == 26788 && 
b[26789] == 26789 && 
b[26790] == 26790 && 
b[26791] == 26791 && 
b[26792] == 26792 && 
b[26793] == 26793 && 
b[26794] == 26794 && 
b[26795] == 26795 && 
b[26796] == 26796 && 
b[26797] == 26797 && 
b[26798] == 26798 && 
b[26799] == 26799 && 
b[26800] == 26800 && 
b[26801] == 26801 && 
b[26802] == 26802 && 
b[26803] == 26803 && 
b[26804] == 26804 && 
b[26805] == 26805 && 
b[26806] == 26806 && 
b[26807] == 26807 && 
b[26808] == 26808 && 
b[26809] == 26809 && 
b[26810] == 26810 && 
b[26811] == 26811 && 
b[26812] == 26812 && 
b[26813] == 26813 && 
b[26814] == 26814 && 
b[26815] == 26815 && 
b[26816] == 26816 && 
b[26817] == 26817 && 
b[26818] == 26818 && 
b[26819] == 26819 && 
b[26820] == 26820 && 
b[26821] == 26821 && 
b[26822] == 26822 && 
b[26823] == 26823 && 
b[26824] == 26824 && 
b[26825] == 26825 && 
b[26826] == 26826 && 
b[26827] == 26827 && 
b[26828] == 26828 && 
b[26829] == 26829 && 
b[26830] == 26830 && 
b[26831] == 26831 && 
b[26832] == 26832 && 
b[26833] == 26833 && 
b[26834] == 26834 && 
b[26835] == 26835 && 
b[26836] == 26836 && 
b[26837] == 26837 && 
b[26838] == 26838 && 
b[26839] == 26839 && 
b[26840] == 26840 && 
b[26841] == 26841 && 
b[26842] == 26842 && 
b[26843] == 26843 && 
b[26844] == 26844 && 
b[26845] == 26845 && 
b[26846] == 26846 && 
b[26847] == 26847 && 
b[26848] == 26848 && 
b[26849] == 26849 && 
b[26850] == 26850 && 
b[26851] == 26851 && 
b[26852] == 26852 && 
b[26853] == 26853 && 
b[26854] == 26854 && 
b[26855] == 26855 && 
b[26856] == 26856 && 
b[26857] == 26857 && 
b[26858] == 26858 && 
b[26859] == 26859 && 
b[26860] == 26860 && 
b[26861] == 26861 && 
b[26862] == 26862 && 
b[26863] == 26863 && 
b[26864] == 26864 && 
b[26865] == 26865 && 
b[26866] == 26866 && 
b[26867] == 26867 && 
b[26868] == 26868 && 
b[26869] == 26869 && 
b[26870] == 26870 && 
b[26871] == 26871 && 
b[26872] == 26872 && 
b[26873] == 26873 && 
b[26874] == 26874 && 
b[26875] == 26875 && 
b[26876] == 26876 && 
b[26877] == 26877 && 
b[26878] == 26878 && 
b[26879] == 26879 && 
b[26880] == 26880 && 
b[26881] == 26881 && 
b[26882] == 26882 && 
b[26883] == 26883 && 
b[26884] == 26884 && 
b[26885] == 26885 && 
b[26886] == 26886 && 
b[26887] == 26887 && 
b[26888] == 26888 && 
b[26889] == 26889 && 
b[26890] == 26890 && 
b[26891] == 26891 && 
b[26892] == 26892 && 
b[26893] == 26893 && 
b[26894] == 26894 && 
b[26895] == 26895 && 
b[26896] == 26896 && 
b[26897] == 26897 && 
b[26898] == 26898 && 
b[26899] == 26899 && 
b[26900] == 26900 && 
b[26901] == 26901 && 
b[26902] == 26902 && 
b[26903] == 26903 && 
b[26904] == 26904 && 
b[26905] == 26905 && 
b[26906] == 26906 && 
b[26907] == 26907 && 
b[26908] == 26908 && 
b[26909] == 26909 && 
b[26910] == 26910 && 
b[26911] == 26911 && 
b[26912] == 26912 && 
b[26913] == 26913 && 
b[26914] == 26914 && 
b[26915] == 26915 && 
b[26916] == 26916 && 
b[26917] == 26917 && 
b[26918] == 26918 && 
b[26919] == 26919 && 
b[26920] == 26920 && 
b[26921] == 26921 && 
b[26922] == 26922 && 
b[26923] == 26923 && 
b[26924] == 26924 && 
b[26925] == 26925 && 
b[26926] == 26926 && 
b[26927] == 26927 && 
b[26928] == 26928 && 
b[26929] == 26929 && 
b[26930] == 26930 && 
b[26931] == 26931 && 
b[26932] == 26932 && 
b[26933] == 26933 && 
b[26934] == 26934 && 
b[26935] == 26935 && 
b[26936] == 26936 && 
b[26937] == 26937 && 
b[26938] == 26938 && 
b[26939] == 26939 && 
b[26940] == 26940 && 
b[26941] == 26941 && 
b[26942] == 26942 && 
b[26943] == 26943 && 
b[26944] == 26944 && 
b[26945] == 26945 && 
b[26946] == 26946 && 
b[26947] == 26947 && 
b[26948] == 26948 && 
b[26949] == 26949 && 
b[26950] == 26950 && 
b[26951] == 26951 && 
b[26952] == 26952 && 
b[26953] == 26953 && 
b[26954] == 26954 && 
b[26955] == 26955 && 
b[26956] == 26956 && 
b[26957] == 26957 && 
b[26958] == 26958 && 
b[26959] == 26959 && 
b[26960] == 26960 && 
b[26961] == 26961 && 
b[26962] == 26962 && 
b[26963] == 26963 && 
b[26964] == 26964 && 
b[26965] == 26965 && 
b[26966] == 26966 && 
b[26967] == 26967 && 
b[26968] == 26968 && 
b[26969] == 26969 && 
b[26970] == 26970 && 
b[26971] == 26971 && 
b[26972] == 26972 && 
b[26973] == 26973 && 
b[26974] == 26974 && 
b[26975] == 26975 && 
b[26976] == 26976 && 
b[26977] == 26977 && 
b[26978] == 26978 && 
b[26979] == 26979 && 
b[26980] == 26980 && 
b[26981] == 26981 && 
b[26982] == 26982 && 
b[26983] == 26983 && 
b[26984] == 26984 && 
b[26985] == 26985 && 
b[26986] == 26986 && 
b[26987] == 26987 && 
b[26988] == 26988 && 
b[26989] == 26989 && 
b[26990] == 26990 && 
b[26991] == 26991 && 
b[26992] == 26992 && 
b[26993] == 26993 && 
b[26994] == 26994 && 
b[26995] == 26995 && 
b[26996] == 26996 && 
b[26997] == 26997 && 
b[26998] == 26998 && 
b[26999] == 26999 && 
b[27000] == 27000 && 
b[27001] == 27001 && 
b[27002] == 27002 && 
b[27003] == 27003 && 
b[27004] == 27004 && 
b[27005] == 27005 && 
b[27006] == 27006 && 
b[27007] == 27007 && 
b[27008] == 27008 && 
b[27009] == 27009 && 
b[27010] == 27010 && 
b[27011] == 27011 && 
b[27012] == 27012 && 
b[27013] == 27013 && 
b[27014] == 27014 && 
b[27015] == 27015 && 
b[27016] == 27016 && 
b[27017] == 27017 && 
b[27018] == 27018 && 
b[27019] == 27019 && 
b[27020] == 27020 && 
b[27021] == 27021 && 
b[27022] == 27022 && 
b[27023] == 27023 && 
b[27024] == 27024 && 
b[27025] == 27025 && 
b[27026] == 27026 && 
b[27027] == 27027 && 
b[27028] == 27028 && 
b[27029] == 27029 && 
b[27030] == 27030 && 
b[27031] == 27031 && 
b[27032] == 27032 && 
b[27033] == 27033 && 
b[27034] == 27034 && 
b[27035] == 27035 && 
b[27036] == 27036 && 
b[27037] == 27037 && 
b[27038] == 27038 && 
b[27039] == 27039 && 
b[27040] == 27040 && 
b[27041] == 27041 && 
b[27042] == 27042 && 
b[27043] == 27043 && 
b[27044] == 27044 && 
b[27045] == 27045 && 
b[27046] == 27046 && 
b[27047] == 27047 && 
b[27048] == 27048 && 
b[27049] == 27049 && 
b[27050] == 27050 && 
b[27051] == 27051 && 
b[27052] == 27052 && 
b[27053] == 27053 && 
b[27054] == 27054 && 
b[27055] == 27055 && 
b[27056] == 27056 && 
b[27057] == 27057 && 
b[27058] == 27058 && 
b[27059] == 27059 && 
b[27060] == 27060 && 
b[27061] == 27061 && 
b[27062] == 27062 && 
b[27063] == 27063 && 
b[27064] == 27064 && 
b[27065] == 27065 && 
b[27066] == 27066 && 
b[27067] == 27067 && 
b[27068] == 27068 && 
b[27069] == 27069 && 
b[27070] == 27070 && 
b[27071] == 27071 && 
b[27072] == 27072 && 
b[27073] == 27073 && 
b[27074] == 27074 && 
b[27075] == 27075 && 
b[27076] == 27076 && 
b[27077] == 27077 && 
b[27078] == 27078 && 
b[27079] == 27079 && 
b[27080] == 27080 && 
b[27081] == 27081 && 
b[27082] == 27082 && 
b[27083] == 27083 && 
b[27084] == 27084 && 
b[27085] == 27085 && 
b[27086] == 27086 && 
b[27087] == 27087 && 
b[27088] == 27088 && 
b[27089] == 27089 && 
b[27090] == 27090 && 
b[27091] == 27091 && 
b[27092] == 27092 && 
b[27093] == 27093 && 
b[27094] == 27094 && 
b[27095] == 27095 && 
b[27096] == 27096 && 
b[27097] == 27097 && 
b[27098] == 27098 && 
b[27099] == 27099 && 
b[27100] == 27100 && 
b[27101] == 27101 && 
b[27102] == 27102 && 
b[27103] == 27103 && 
b[27104] == 27104 && 
b[27105] == 27105 && 
b[27106] == 27106 && 
b[27107] == 27107 && 
b[27108] == 27108 && 
b[27109] == 27109 && 
b[27110] == 27110 && 
b[27111] == 27111 && 
b[27112] == 27112 && 
b[27113] == 27113 && 
b[27114] == 27114 && 
b[27115] == 27115 && 
b[27116] == 27116 && 
b[27117] == 27117 && 
b[27118] == 27118 && 
b[27119] == 27119 && 
b[27120] == 27120 && 
b[27121] == 27121 && 
b[27122] == 27122 && 
b[27123] == 27123 && 
b[27124] == 27124 && 
b[27125] == 27125 && 
b[27126] == 27126 && 
b[27127] == 27127 && 
b[27128] == 27128 && 
b[27129] == 27129 && 
b[27130] == 27130 && 
b[27131] == 27131 && 
b[27132] == 27132 && 
b[27133] == 27133 && 
b[27134] == 27134 && 
b[27135] == 27135 && 
b[27136] == 27136 && 
b[27137] == 27137 && 
b[27138] == 27138 && 
b[27139] == 27139 && 
b[27140] == 27140 && 
b[27141] == 27141 && 
b[27142] == 27142 && 
b[27143] == 27143 && 
b[27144] == 27144 && 
b[27145] == 27145 && 
b[27146] == 27146 && 
b[27147] == 27147 && 
b[27148] == 27148 && 
b[27149] == 27149 && 
b[27150] == 27150 && 
b[27151] == 27151 && 
b[27152] == 27152 && 
b[27153] == 27153 && 
b[27154] == 27154 && 
b[27155] == 27155 && 
b[27156] == 27156 && 
b[27157] == 27157 && 
b[27158] == 27158 && 
b[27159] == 27159 && 
b[27160] == 27160 && 
b[27161] == 27161 && 
b[27162] == 27162 && 
b[27163] == 27163 && 
b[27164] == 27164 && 
b[27165] == 27165 && 
b[27166] == 27166 && 
b[27167] == 27167 && 
b[27168] == 27168 && 
b[27169] == 27169 && 
b[27170] == 27170 && 
b[27171] == 27171 && 
b[27172] == 27172 && 
b[27173] == 27173 && 
b[27174] == 27174 && 
b[27175] == 27175 && 
b[27176] == 27176 && 
b[27177] == 27177 && 
b[27178] == 27178 && 
b[27179] == 27179 && 
b[27180] == 27180 && 
b[27181] == 27181 && 
b[27182] == 27182 && 
b[27183] == 27183 && 
b[27184] == 27184 && 
b[27185] == 27185 && 
b[27186] == 27186 && 
b[27187] == 27187 && 
b[27188] == 27188 && 
b[27189] == 27189 && 
b[27190] == 27190 && 
b[27191] == 27191 && 
b[27192] == 27192 && 
b[27193] == 27193 && 
b[27194] == 27194 && 
b[27195] == 27195 && 
b[27196] == 27196 && 
b[27197] == 27197 && 
b[27198] == 27198 && 
b[27199] == 27199 && 
b[27200] == 27200 && 
b[27201] == 27201 && 
b[27202] == 27202 && 
b[27203] == 27203 && 
b[27204] == 27204 && 
b[27205] == 27205 && 
b[27206] == 27206 && 
b[27207] == 27207 && 
b[27208] == 27208 && 
b[27209] == 27209 && 
b[27210] == 27210 && 
b[27211] == 27211 && 
b[27212] == 27212 && 
b[27213] == 27213 && 
b[27214] == 27214 && 
b[27215] == 27215 && 
b[27216] == 27216 && 
b[27217] == 27217 && 
b[27218] == 27218 && 
b[27219] == 27219 && 
b[27220] == 27220 && 
b[27221] == 27221 && 
b[27222] == 27222 && 
b[27223] == 27223 && 
b[27224] == 27224 && 
b[27225] == 27225 && 
b[27226] == 27226 && 
b[27227] == 27227 && 
b[27228] == 27228 && 
b[27229] == 27229 && 
b[27230] == 27230 && 
b[27231] == 27231 && 
b[27232] == 27232 && 
b[27233] == 27233 && 
b[27234] == 27234 && 
b[27235] == 27235 && 
b[27236] == 27236 && 
b[27237] == 27237 && 
b[27238] == 27238 && 
b[27239] == 27239 && 
b[27240] == 27240 && 
b[27241] == 27241 && 
b[27242] == 27242 && 
b[27243] == 27243 && 
b[27244] == 27244 && 
b[27245] == 27245 && 
b[27246] == 27246 && 
b[27247] == 27247 && 
b[27248] == 27248 && 
b[27249] == 27249 && 
b[27250] == 27250 && 
b[27251] == 27251 && 
b[27252] == 27252 && 
b[27253] == 27253 && 
b[27254] == 27254 && 
b[27255] == 27255 && 
b[27256] == 27256 && 
b[27257] == 27257 && 
b[27258] == 27258 && 
b[27259] == 27259 && 
b[27260] == 27260 && 
b[27261] == 27261 && 
b[27262] == 27262 && 
b[27263] == 27263 && 
b[27264] == 27264 && 
b[27265] == 27265 && 
b[27266] == 27266 && 
b[27267] == 27267 && 
b[27268] == 27268 && 
b[27269] == 27269 && 
b[27270] == 27270 && 
b[27271] == 27271 && 
b[27272] == 27272 && 
b[27273] == 27273 && 
b[27274] == 27274 && 
b[27275] == 27275 && 
b[27276] == 27276 && 
b[27277] == 27277 && 
b[27278] == 27278 && 
b[27279] == 27279 && 
b[27280] == 27280 && 
b[27281] == 27281 && 
b[27282] == 27282 && 
b[27283] == 27283 && 
b[27284] == 27284 && 
b[27285] == 27285 && 
b[27286] == 27286 && 
b[27287] == 27287 && 
b[27288] == 27288 && 
b[27289] == 27289 && 
b[27290] == 27290 && 
b[27291] == 27291 && 
b[27292] == 27292 && 
b[27293] == 27293 && 
b[27294] == 27294 && 
b[27295] == 27295 && 
b[27296] == 27296 && 
b[27297] == 27297 && 
b[27298] == 27298 && 
b[27299] == 27299 && 
b[27300] == 27300 && 
b[27301] == 27301 && 
b[27302] == 27302 && 
b[27303] == 27303 && 
b[27304] == 27304 && 
b[27305] == 27305 && 
b[27306] == 27306 && 
b[27307] == 27307 && 
b[27308] == 27308 && 
b[27309] == 27309 && 
b[27310] == 27310 && 
b[27311] == 27311 && 
b[27312] == 27312 && 
b[27313] == 27313 && 
b[27314] == 27314 && 
b[27315] == 27315 && 
b[27316] == 27316 && 
b[27317] == 27317 && 
b[27318] == 27318 && 
b[27319] == 27319 && 
b[27320] == 27320 && 
b[27321] == 27321 && 
b[27322] == 27322 && 
b[27323] == 27323 && 
b[27324] == 27324 && 
b[27325] == 27325 && 
b[27326] == 27326 && 
b[27327] == 27327 && 
b[27328] == 27328 && 
b[27329] == 27329 && 
b[27330] == 27330 && 
b[27331] == 27331 && 
b[27332] == 27332 && 
b[27333] == 27333 && 
b[27334] == 27334 && 
b[27335] == 27335 && 
b[27336] == 27336 && 
b[27337] == 27337 && 
b[27338] == 27338 && 
b[27339] == 27339 && 
b[27340] == 27340 && 
b[27341] == 27341 && 
b[27342] == 27342 && 
b[27343] == 27343 && 
b[27344] == 27344 && 
b[27345] == 27345 && 
b[27346] == 27346 && 
b[27347] == 27347 && 
b[27348] == 27348 && 
b[27349] == 27349 && 
b[27350] == 27350 && 
b[27351] == 27351 && 
b[27352] == 27352 && 
b[27353] == 27353 && 
b[27354] == 27354 && 
b[27355] == 27355 && 
b[27356] == 27356 && 
b[27357] == 27357 && 
b[27358] == 27358 && 
b[27359] == 27359 && 
b[27360] == 27360 && 
b[27361] == 27361 && 
b[27362] == 27362 && 
b[27363] == 27363 && 
b[27364] == 27364 && 
b[27365] == 27365 && 
b[27366] == 27366 && 
b[27367] == 27367 && 
b[27368] == 27368 && 
b[27369] == 27369 && 
b[27370] == 27370 && 
b[27371] == 27371 && 
b[27372] == 27372 && 
b[27373] == 27373 && 
b[27374] == 27374 && 
b[27375] == 27375 && 
b[27376] == 27376 && 
b[27377] == 27377 && 
b[27378] == 27378 && 
b[27379] == 27379 && 
b[27380] == 27380 && 
b[27381] == 27381 && 
b[27382] == 27382 && 
b[27383] == 27383 && 
b[27384] == 27384 && 
b[27385] == 27385 && 
b[27386] == 27386 && 
b[27387] == 27387 && 
b[27388] == 27388 && 
b[27389] == 27389 && 
b[27390] == 27390 && 
b[27391] == 27391 && 
b[27392] == 27392 && 
b[27393] == 27393 && 
b[27394] == 27394 && 
b[27395] == 27395 && 
b[27396] == 27396 && 
b[27397] == 27397 && 
b[27398] == 27398 && 
b[27399] == 27399 && 
b[27400] == 27400 && 
b[27401] == 27401 && 
b[27402] == 27402 && 
b[27403] == 27403 && 
b[27404] == 27404 && 
b[27405] == 27405 && 
b[27406] == 27406 && 
b[27407] == 27407 && 
b[27408] == 27408 && 
b[27409] == 27409 && 
b[27410] == 27410 && 
b[27411] == 27411 && 
b[27412] == 27412 && 
b[27413] == 27413 && 
b[27414] == 27414 && 
b[27415] == 27415 && 
b[27416] == 27416 && 
b[27417] == 27417 && 
b[27418] == 27418 && 
b[27419] == 27419 && 
b[27420] == 27420 && 
b[27421] == 27421 && 
b[27422] == 27422 && 
b[27423] == 27423 && 
b[27424] == 27424 && 
b[27425] == 27425 && 
b[27426] == 27426 && 
b[27427] == 27427 && 
b[27428] == 27428 && 
b[27429] == 27429 && 
b[27430] == 27430 && 
b[27431] == 27431 && 
b[27432] == 27432 && 
b[27433] == 27433 && 
b[27434] == 27434 && 
b[27435] == 27435 && 
b[27436] == 27436 && 
b[27437] == 27437 && 
b[27438] == 27438 && 
b[27439] == 27439 && 
b[27440] == 27440 && 
b[27441] == 27441 && 
b[27442] == 27442 && 
b[27443] == 27443 && 
b[27444] == 27444 && 
b[27445] == 27445 && 
b[27446] == 27446 && 
b[27447] == 27447 && 
b[27448] == 27448 && 
b[27449] == 27449 && 
b[27450] == 27450 && 
b[27451] == 27451 && 
b[27452] == 27452 && 
b[27453] == 27453 && 
b[27454] == 27454 && 
b[27455] == 27455 && 
b[27456] == 27456 && 
b[27457] == 27457 && 
b[27458] == 27458 && 
b[27459] == 27459 && 
b[27460] == 27460 && 
b[27461] == 27461 && 
b[27462] == 27462 && 
b[27463] == 27463 && 
b[27464] == 27464 && 
b[27465] == 27465 && 
b[27466] == 27466 && 
b[27467] == 27467 && 
b[27468] == 27468 && 
b[27469] == 27469 && 
b[27470] == 27470 && 
b[27471] == 27471 && 
b[27472] == 27472 && 
b[27473] == 27473 && 
b[27474] == 27474 && 
b[27475] == 27475 && 
b[27476] == 27476 && 
b[27477] == 27477 && 
b[27478] == 27478 && 
b[27479] == 27479 && 
b[27480] == 27480 && 
b[27481] == 27481 && 
b[27482] == 27482 && 
b[27483] == 27483 && 
b[27484] == 27484 && 
b[27485] == 27485 && 
b[27486] == 27486 && 
b[27487] == 27487 && 
b[27488] == 27488 && 
b[27489] == 27489 && 
b[27490] == 27490 && 
b[27491] == 27491 && 
b[27492] == 27492 && 
b[27493] == 27493 && 
b[27494] == 27494 && 
b[27495] == 27495 && 
b[27496] == 27496 && 
b[27497] == 27497 && 
b[27498] == 27498 && 
b[27499] == 27499 && 
b[27500] == 27500 && 
b[27501] == 27501 && 
b[27502] == 27502 && 
b[27503] == 27503 && 
b[27504] == 27504 && 
b[27505] == 27505 && 
b[27506] == 27506 && 
b[27507] == 27507 && 
b[27508] == 27508 && 
b[27509] == 27509 && 
b[27510] == 27510 && 
b[27511] == 27511 && 
b[27512] == 27512 && 
b[27513] == 27513 && 
b[27514] == 27514 && 
b[27515] == 27515 && 
b[27516] == 27516 && 
b[27517] == 27517 && 
b[27518] == 27518 && 
b[27519] == 27519 && 
b[27520] == 27520 && 
b[27521] == 27521 && 
b[27522] == 27522 && 
b[27523] == 27523 && 
b[27524] == 27524 && 
b[27525] == 27525 && 
b[27526] == 27526 && 
b[27527] == 27527 && 
b[27528] == 27528 && 
b[27529] == 27529 && 
b[27530] == 27530 && 
b[27531] == 27531 && 
b[27532] == 27532 && 
b[27533] == 27533 && 
b[27534] == 27534 && 
b[27535] == 27535 && 
b[27536] == 27536 && 
b[27537] == 27537 && 
b[27538] == 27538 && 
b[27539] == 27539 && 
b[27540] == 27540 && 
b[27541] == 27541 && 
b[27542] == 27542 && 
b[27543] == 27543 && 
b[27544] == 27544 && 
b[27545] == 27545 && 
b[27546] == 27546 && 
b[27547] == 27547 && 
b[27548] == 27548 && 
b[27549] == 27549 && 
b[27550] == 27550 && 
b[27551] == 27551 && 
b[27552] == 27552 && 
b[27553] == 27553 && 
b[27554] == 27554 && 
b[27555] == 27555 && 
b[27556] == 27556 && 
b[27557] == 27557 && 
b[27558] == 27558 && 
b[27559] == 27559 && 
b[27560] == 27560 && 
b[27561] == 27561 && 
b[27562] == 27562 && 
b[27563] == 27563 && 
b[27564] == 27564 && 
b[27565] == 27565 && 
b[27566] == 27566 && 
b[27567] == 27567 && 
b[27568] == 27568 && 
b[27569] == 27569 && 
b[27570] == 27570 && 
b[27571] == 27571 && 
b[27572] == 27572 && 
b[27573] == 27573 && 
b[27574] == 27574 && 
b[27575] == 27575 && 
b[27576] == 27576 && 
b[27577] == 27577 && 
b[27578] == 27578 && 
b[27579] == 27579 && 
b[27580] == 27580 && 
b[27581] == 27581 && 
b[27582] == 27582 && 
b[27583] == 27583 && 
b[27584] == 27584 && 
b[27585] == 27585 && 
b[27586] == 27586 && 
b[27587] == 27587 && 
b[27588] == 27588 && 
b[27589] == 27589 && 
b[27590] == 27590 && 
b[27591] == 27591 && 
b[27592] == 27592 && 
b[27593] == 27593 && 
b[27594] == 27594 && 
b[27595] == 27595 && 
b[27596] == 27596 && 
b[27597] == 27597 && 
b[27598] == 27598 && 
b[27599] == 27599 && 
b[27600] == 27600 && 
b[27601] == 27601 && 
b[27602] == 27602 && 
b[27603] == 27603 && 
b[27604] == 27604 && 
b[27605] == 27605 && 
b[27606] == 27606 && 
b[27607] == 27607 && 
b[27608] == 27608 && 
b[27609] == 27609 && 
b[27610] == 27610 && 
b[27611] == 27611 && 
b[27612] == 27612 && 
b[27613] == 27613 && 
b[27614] == 27614 && 
b[27615] == 27615 && 
b[27616] == 27616 && 
b[27617] == 27617 && 
b[27618] == 27618 && 
b[27619] == 27619 && 
b[27620] == 27620 && 
b[27621] == 27621 && 
b[27622] == 27622 && 
b[27623] == 27623 && 
b[27624] == 27624 && 
b[27625] == 27625 && 
b[27626] == 27626 && 
b[27627] == 27627 && 
b[27628] == 27628 && 
b[27629] == 27629 && 
b[27630] == 27630 && 
b[27631] == 27631 && 
b[27632] == 27632 && 
b[27633] == 27633 && 
b[27634] == 27634 && 
b[27635] == 27635 && 
b[27636] == 27636 && 
b[27637] == 27637 && 
b[27638] == 27638 && 
b[27639] == 27639 && 
b[27640] == 27640 && 
b[27641] == 27641 && 
b[27642] == 27642 && 
b[27643] == 27643 && 
b[27644] == 27644 && 
b[27645] == 27645 && 
b[27646] == 27646 && 
b[27647] == 27647 && 
b[27648] == 27648 && 
b[27649] == 27649 && 
b[27650] == 27650 && 
b[27651] == 27651 && 
b[27652] == 27652 && 
b[27653] == 27653 && 
b[27654] == 27654 && 
b[27655] == 27655 && 
b[27656] == 27656 && 
b[27657] == 27657 && 
b[27658] == 27658 && 
b[27659] == 27659 && 
b[27660] == 27660 && 
b[27661] == 27661 && 
b[27662] == 27662 && 
b[27663] == 27663 && 
b[27664] == 27664 && 
b[27665] == 27665 && 
b[27666] == 27666 && 
b[27667] == 27667 && 
b[27668] == 27668 && 
b[27669] == 27669 && 
b[27670] == 27670 && 
b[27671] == 27671 && 
b[27672] == 27672 && 
b[27673] == 27673 && 
b[27674] == 27674 && 
b[27675] == 27675 && 
b[27676] == 27676 && 
b[27677] == 27677 && 
b[27678] == 27678 && 
b[27679] == 27679 && 
b[27680] == 27680 && 
b[27681] == 27681 && 
b[27682] == 27682 && 
b[27683] == 27683 && 
b[27684] == 27684 && 
b[27685] == 27685 && 
b[27686] == 27686 && 
b[27687] == 27687 && 
b[27688] == 27688 && 
b[27689] == 27689 && 
b[27690] == 27690 && 
b[27691] == 27691 && 
b[27692] == 27692 && 
b[27693] == 27693 && 
b[27694] == 27694 && 
b[27695] == 27695 && 
b[27696] == 27696 && 
b[27697] == 27697 && 
b[27698] == 27698 && 
b[27699] == 27699 && 
b[27700] == 27700 && 
b[27701] == 27701 && 
b[27702] == 27702 && 
b[27703] == 27703 && 
b[27704] == 27704 && 
b[27705] == 27705 && 
b[27706] == 27706 && 
b[27707] == 27707 && 
b[27708] == 27708 && 
b[27709] == 27709 && 
b[27710] == 27710 && 
b[27711] == 27711 && 
b[27712] == 27712 && 
b[27713] == 27713 && 
b[27714] == 27714 && 
b[27715] == 27715 && 
b[27716] == 27716 && 
b[27717] == 27717 && 
b[27718] == 27718 && 
b[27719] == 27719 && 
b[27720] == 27720 && 
b[27721] == 27721 && 
b[27722] == 27722 && 
b[27723] == 27723 && 
b[27724] == 27724 && 
b[27725] == 27725 && 
b[27726] == 27726 && 
b[27727] == 27727 && 
b[27728] == 27728 && 
b[27729] == 27729 && 
b[27730] == 27730 && 
b[27731] == 27731 && 
b[27732] == 27732 && 
b[27733] == 27733 && 
b[27734] == 27734 && 
b[27735] == 27735 && 
b[27736] == 27736 && 
b[27737] == 27737 && 
b[27738] == 27738 && 
b[27739] == 27739 && 
b[27740] == 27740 && 
b[27741] == 27741 && 
b[27742] == 27742 && 
b[27743] == 27743 && 
b[27744] == 27744 && 
b[27745] == 27745 && 
b[27746] == 27746 && 
b[27747] == 27747 && 
b[27748] == 27748 && 
b[27749] == 27749 && 
b[27750] == 27750 && 
b[27751] == 27751 && 
b[27752] == 27752 && 
b[27753] == 27753 && 
b[27754] == 27754 && 
b[27755] == 27755 && 
b[27756] == 27756 && 
b[27757] == 27757 && 
b[27758] == 27758 && 
b[27759] == 27759 && 
b[27760] == 27760 && 
b[27761] == 27761 && 
b[27762] == 27762 && 
b[27763] == 27763 && 
b[27764] == 27764 && 
b[27765] == 27765 && 
b[27766] == 27766 && 
b[27767] == 27767 && 
b[27768] == 27768 && 
b[27769] == 27769 && 
b[27770] == 27770 && 
b[27771] == 27771 && 
b[27772] == 27772 && 
b[27773] == 27773 && 
b[27774] == 27774 && 
b[27775] == 27775 && 
b[27776] == 27776 && 
b[27777] == 27777 && 
b[27778] == 27778 && 
b[27779] == 27779 && 
b[27780] == 27780 && 
b[27781] == 27781 && 
b[27782] == 27782 && 
b[27783] == 27783 && 
b[27784] == 27784 && 
b[27785] == 27785 && 
b[27786] == 27786 && 
b[27787] == 27787 && 
b[27788] == 27788 && 
b[27789] == 27789 && 
b[27790] == 27790 && 
b[27791] == 27791 && 
b[27792] == 27792 && 
b[27793] == 27793 && 
b[27794] == 27794 && 
b[27795] == 27795 && 
b[27796] == 27796 && 
b[27797] == 27797 && 
b[27798] == 27798 && 
b[27799] == 27799 && 
b[27800] == 27800 && 
b[27801] == 27801 && 
b[27802] == 27802 && 
b[27803] == 27803 && 
b[27804] == 27804 && 
b[27805] == 27805 && 
b[27806] == 27806 && 
b[27807] == 27807 && 
b[27808] == 27808 && 
b[27809] == 27809 && 
b[27810] == 27810 && 
b[27811] == 27811 && 
b[27812] == 27812 && 
b[27813] == 27813 && 
b[27814] == 27814 && 
b[27815] == 27815 && 
b[27816] == 27816 && 
b[27817] == 27817 && 
b[27818] == 27818 && 
b[27819] == 27819 && 
b[27820] == 27820 && 
b[27821] == 27821 && 
b[27822] == 27822 && 
b[27823] == 27823 && 
b[27824] == 27824 && 
b[27825] == 27825 && 
b[27826] == 27826 && 
b[27827] == 27827 && 
b[27828] == 27828 && 
b[27829] == 27829 && 
b[27830] == 27830 && 
b[27831] == 27831 && 
b[27832] == 27832 && 
b[27833] == 27833 && 
b[27834] == 27834 && 
b[27835] == 27835 && 
b[27836] == 27836 && 
b[27837] == 27837 && 
b[27838] == 27838 && 
b[27839] == 27839 && 
b[27840] == 27840 && 
b[27841] == 27841 && 
b[27842] == 27842 && 
b[27843] == 27843 && 
b[27844] == 27844 && 
b[27845] == 27845 && 
b[27846] == 27846 && 
b[27847] == 27847 && 
b[27848] == 27848 && 
b[27849] == 27849 && 
b[27850] == 27850 && 
b[27851] == 27851 && 
b[27852] == 27852 && 
b[27853] == 27853 && 
b[27854] == 27854 && 
b[27855] == 27855 && 
b[27856] == 27856 && 
b[27857] == 27857 && 
b[27858] == 27858 && 
b[27859] == 27859 && 
b[27860] == 27860 && 
b[27861] == 27861 && 
b[27862] == 27862 && 
b[27863] == 27863 && 
b[27864] == 27864 && 
b[27865] == 27865 && 
b[27866] == 27866 && 
b[27867] == 27867 && 
b[27868] == 27868 && 
b[27869] == 27869 && 
b[27870] == 27870 && 
b[27871] == 27871 && 
b[27872] == 27872 && 
b[27873] == 27873 && 
b[27874] == 27874 && 
b[27875] == 27875 && 
b[27876] == 27876 && 
b[27877] == 27877 && 
b[27878] == 27878 && 
b[27879] == 27879 && 
b[27880] == 27880 && 
b[27881] == 27881 && 
b[27882] == 27882 && 
b[27883] == 27883 && 
b[27884] == 27884 && 
b[27885] == 27885 && 
b[27886] == 27886 && 
b[27887] == 27887 && 
b[27888] == 27888 && 
b[27889] == 27889 && 
b[27890] == 27890 && 
b[27891] == 27891 && 
b[27892] == 27892 && 
b[27893] == 27893 && 
b[27894] == 27894 && 
b[27895] == 27895 && 
b[27896] == 27896 && 
b[27897] == 27897 && 
b[27898] == 27898 && 
b[27899] == 27899 && 
b[27900] == 27900 && 
b[27901] == 27901 && 
b[27902] == 27902 && 
b[27903] == 27903 && 
b[27904] == 27904 && 
b[27905] == 27905 && 
b[27906] == 27906 && 
b[27907] == 27907 && 
b[27908] == 27908 && 
b[27909] == 27909 && 
b[27910] == 27910 && 
b[27911] == 27911 && 
b[27912] == 27912 && 
b[27913] == 27913 && 
b[27914] == 27914 && 
b[27915] == 27915 && 
b[27916] == 27916 && 
b[27917] == 27917 && 
b[27918] == 27918 && 
b[27919] == 27919 && 
b[27920] == 27920 && 
b[27921] == 27921 && 
b[27922] == 27922 && 
b[27923] == 27923 && 
b[27924] == 27924 && 
b[27925] == 27925 && 
b[27926] == 27926 && 
b[27927] == 27927 && 
b[27928] == 27928 && 
b[27929] == 27929 && 
b[27930] == 27930 && 
b[27931] == 27931 && 
b[27932] == 27932 && 
b[27933] == 27933 && 
b[27934] == 27934 && 
b[27935] == 27935 && 
b[27936] == 27936 && 
b[27937] == 27937 && 
b[27938] == 27938 && 
b[27939] == 27939 && 
b[27940] == 27940 && 
b[27941] == 27941 && 
b[27942] == 27942 && 
b[27943] == 27943 && 
b[27944] == 27944 && 
b[27945] == 27945 && 
b[27946] == 27946 && 
b[27947] == 27947 && 
b[27948] == 27948 && 
b[27949] == 27949 && 
b[27950] == 27950 && 
b[27951] == 27951 && 
b[27952] == 27952 && 
b[27953] == 27953 && 
b[27954] == 27954 && 
b[27955] == 27955 && 
b[27956] == 27956 && 
b[27957] == 27957 && 
b[27958] == 27958 && 
b[27959] == 27959 && 
b[27960] == 27960 && 
b[27961] == 27961 && 
b[27962] == 27962 && 
b[27963] == 27963 && 
b[27964] == 27964 && 
b[27965] == 27965 && 
b[27966] == 27966 && 
b[27967] == 27967 && 
b[27968] == 27968 && 
b[27969] == 27969 && 
b[27970] == 27970 && 
b[27971] == 27971 && 
b[27972] == 27972 && 
b[27973] == 27973 && 
b[27974] == 27974 && 
b[27975] == 27975 && 
b[27976] == 27976 && 
b[27977] == 27977 && 
b[27978] == 27978 && 
b[27979] == 27979 && 
b[27980] == 27980 && 
b[27981] == 27981 && 
b[27982] == 27982 && 
b[27983] == 27983 && 
b[27984] == 27984 && 
b[27985] == 27985 && 
b[27986] == 27986 && 
b[27987] == 27987 && 
b[27988] == 27988 && 
b[27989] == 27989 && 
b[27990] == 27990 && 
b[27991] == 27991 && 
b[27992] == 27992 && 
b[27993] == 27993 && 
b[27994] == 27994 && 
b[27995] == 27995 && 
b[27996] == 27996 && 
b[27997] == 27997 && 
b[27998] == 27998 && 
b[27999] == 27999 && 
b[28000] == 28000 && 
b[28001] == 28001 && 
b[28002] == 28002 && 
b[28003] == 28003 && 
b[28004] == 28004 && 
b[28005] == 28005 && 
b[28006] == 28006 && 
b[28007] == 28007 && 
b[28008] == 28008 && 
b[28009] == 28009 && 
b[28010] == 28010 && 
b[28011] == 28011 && 
b[28012] == 28012 && 
b[28013] == 28013 && 
b[28014] == 28014 && 
b[28015] == 28015 && 
b[28016] == 28016 && 
b[28017] == 28017 && 
b[28018] == 28018 && 
b[28019] == 28019 && 
b[28020] == 28020 && 
b[28021] == 28021 && 
b[28022] == 28022 && 
b[28023] == 28023 && 
b[28024] == 28024 && 
b[28025] == 28025 && 
b[28026] == 28026 && 
b[28027] == 28027 && 
b[28028] == 28028 && 
b[28029] == 28029 && 
b[28030] == 28030 && 
b[28031] == 28031 && 
b[28032] == 28032 && 
b[28033] == 28033 && 
b[28034] == 28034 && 
b[28035] == 28035 && 
b[28036] == 28036 && 
b[28037] == 28037 && 
b[28038] == 28038 && 
b[28039] == 28039 && 
b[28040] == 28040 && 
b[28041] == 28041 && 
b[28042] == 28042 && 
b[28043] == 28043 && 
b[28044] == 28044 && 
b[28045] == 28045 && 
b[28046] == 28046 && 
b[28047] == 28047 && 
b[28048] == 28048 && 
b[28049] == 28049 && 
b[28050] == 28050 && 
b[28051] == 28051 && 
b[28052] == 28052 && 
b[28053] == 28053 && 
b[28054] == 28054 && 
b[28055] == 28055 && 
b[28056] == 28056 && 
b[28057] == 28057 && 
b[28058] == 28058 && 
b[28059] == 28059 && 
b[28060] == 28060 && 
b[28061] == 28061 && 
b[28062] == 28062 && 
b[28063] == 28063 && 
b[28064] == 28064 && 
b[28065] == 28065 && 
b[28066] == 28066 && 
b[28067] == 28067 && 
b[28068] == 28068 && 
b[28069] == 28069 && 
b[28070] == 28070 && 
b[28071] == 28071 && 
b[28072] == 28072 && 
b[28073] == 28073 && 
b[28074] == 28074 && 
b[28075] == 28075 && 
b[28076] == 28076 && 
b[28077] == 28077 && 
b[28078] == 28078 && 
b[28079] == 28079 && 
b[28080] == 28080 && 
b[28081] == 28081 && 
b[28082] == 28082 && 
b[28083] == 28083 && 
b[28084] == 28084 && 
b[28085] == 28085 && 
b[28086] == 28086 && 
b[28087] == 28087 && 
b[28088] == 28088 && 
b[28089] == 28089 && 
b[28090] == 28090 && 
b[28091] == 28091 && 
b[28092] == 28092 && 
b[28093] == 28093 && 
b[28094] == 28094 && 
b[28095] == 28095 && 
b[28096] == 28096 && 
b[28097] == 28097 && 
b[28098] == 28098 && 
b[28099] == 28099 && 
b[28100] == 28100 && 
b[28101] == 28101 && 
b[28102] == 28102 && 
b[28103] == 28103 && 
b[28104] == 28104 && 
b[28105] == 28105 && 
b[28106] == 28106 && 
b[28107] == 28107 && 
b[28108] == 28108 && 
b[28109] == 28109 && 
b[28110] == 28110 && 
b[28111] == 28111 && 
b[28112] == 28112 && 
b[28113] == 28113 && 
b[28114] == 28114 && 
b[28115] == 28115 && 
b[28116] == 28116 && 
b[28117] == 28117 && 
b[28118] == 28118 && 
b[28119] == 28119 && 
b[28120] == 28120 && 
b[28121] == 28121 && 
b[28122] == 28122 && 
b[28123] == 28123 && 
b[28124] == 28124 && 
b[28125] == 28125 && 
b[28126] == 28126 && 
b[28127] == 28127 && 
b[28128] == 28128 && 
b[28129] == 28129 && 
b[28130] == 28130 && 
b[28131] == 28131 && 
b[28132] == 28132 && 
b[28133] == 28133 && 
b[28134] == 28134 && 
b[28135] == 28135 && 
b[28136] == 28136 && 
b[28137] == 28137 && 
b[28138] == 28138 && 
b[28139] == 28139 && 
b[28140] == 28140 && 
b[28141] == 28141 && 
b[28142] == 28142 && 
b[28143] == 28143 && 
b[28144] == 28144 && 
b[28145] == 28145 && 
b[28146] == 28146 && 
b[28147] == 28147 && 
b[28148] == 28148 && 
b[28149] == 28149 && 
b[28150] == 28150 && 
b[28151] == 28151 && 
b[28152] == 28152 && 
b[28153] == 28153 && 
b[28154] == 28154 && 
b[28155] == 28155 && 
b[28156] == 28156 && 
b[28157] == 28157 && 
b[28158] == 28158 && 
b[28159] == 28159 && 
b[28160] == 28160 && 
b[28161] == 28161 && 
b[28162] == 28162 && 
b[28163] == 28163 && 
b[28164] == 28164 && 
b[28165] == 28165 && 
b[28166] == 28166 && 
b[28167] == 28167 && 
b[28168] == 28168 && 
b[28169] == 28169 && 
b[28170] == 28170 && 
b[28171] == 28171 && 
b[28172] == 28172 && 
b[28173] == 28173 && 
b[28174] == 28174 && 
b[28175] == 28175 && 
b[28176] == 28176 && 
b[28177] == 28177 && 
b[28178] == 28178 && 
b[28179] == 28179 && 
b[28180] == 28180 && 
b[28181] == 28181 && 
b[28182] == 28182 && 
b[28183] == 28183 && 
b[28184] == 28184 && 
b[28185] == 28185 && 
b[28186] == 28186 && 
b[28187] == 28187 && 
b[28188] == 28188 && 
b[28189] == 28189 && 
b[28190] == 28190 && 
b[28191] == 28191 && 
b[28192] == 28192 && 
b[28193] == 28193 && 
b[28194] == 28194 && 
b[28195] == 28195 && 
b[28196] == 28196 && 
b[28197] == 28197 && 
b[28198] == 28198 && 
b[28199] == 28199 && 
b[28200] == 28200 && 
b[28201] == 28201 && 
b[28202] == 28202 && 
b[28203] == 28203 && 
b[28204] == 28204 && 
b[28205] == 28205 && 
b[28206] == 28206 && 
b[28207] == 28207 && 
b[28208] == 28208 && 
b[28209] == 28209 && 
b[28210] == 28210 && 
b[28211] == 28211 && 
b[28212] == 28212 && 
b[28213] == 28213 && 
b[28214] == 28214 && 
b[28215] == 28215 && 
b[28216] == 28216 && 
b[28217] == 28217 && 
b[28218] == 28218 && 
b[28219] == 28219 && 
b[28220] == 28220 && 
b[28221] == 28221 && 
b[28222] == 28222 && 
b[28223] == 28223 && 
b[28224] == 28224 && 
b[28225] == 28225 && 
b[28226] == 28226 && 
b[28227] == 28227 && 
b[28228] == 28228 && 
b[28229] == 28229 && 
b[28230] == 28230 && 
b[28231] == 28231 && 
b[28232] == 28232 && 
b[28233] == 28233 && 
b[28234] == 28234 && 
b[28235] == 28235 && 
b[28236] == 28236 && 
b[28237] == 28237 && 
b[28238] == 28238 && 
b[28239] == 28239 && 
b[28240] == 28240 && 
b[28241] == 28241 && 
b[28242] == 28242 && 
b[28243] == 28243 && 
b[28244] == 28244 && 
b[28245] == 28245 && 
b[28246] == 28246 && 
b[28247] == 28247 && 
b[28248] == 28248 && 
b[28249] == 28249 && 
b[28250] == 28250 && 
b[28251] == 28251 && 
b[28252] == 28252 && 
b[28253] == 28253 && 
b[28254] == 28254 && 
b[28255] == 28255 && 
b[28256] == 28256 && 
b[28257] == 28257 && 
b[28258] == 28258 && 
b[28259] == 28259 && 
b[28260] == 28260 && 
b[28261] == 28261 && 
b[28262] == 28262 && 
b[28263] == 28263 && 
b[28264] == 28264 && 
b[28265] == 28265 && 
b[28266] == 28266 && 
b[28267] == 28267 && 
b[28268] == 28268 && 
b[28269] == 28269 && 
b[28270] == 28270 && 
b[28271] == 28271 && 
b[28272] == 28272 && 
b[28273] == 28273 && 
b[28274] == 28274 && 
b[28275] == 28275 && 
b[28276] == 28276 && 
b[28277] == 28277 && 
b[28278] == 28278 && 
b[28279] == 28279 && 
b[28280] == 28280 && 
b[28281] == 28281 && 
b[28282] == 28282 && 
b[28283] == 28283 && 
b[28284] == 28284 && 
b[28285] == 28285 && 
b[28286] == 28286 && 
b[28287] == 28287 && 
b[28288] == 28288 && 
b[28289] == 28289 && 
b[28290] == 28290 && 
b[28291] == 28291 && 
b[28292] == 28292 && 
b[28293] == 28293 && 
b[28294] == 28294 && 
b[28295] == 28295 && 
b[28296] == 28296 && 
b[28297] == 28297 && 
b[28298] == 28298 && 
b[28299] == 28299 && 
b[28300] == 28300 && 
b[28301] == 28301 && 
b[28302] == 28302 && 
b[28303] == 28303 && 
b[28304] == 28304 && 
b[28305] == 28305 && 
b[28306] == 28306 && 
b[28307] == 28307 && 
b[28308] == 28308 && 
b[28309] == 28309 && 
b[28310] == 28310 && 
b[28311] == 28311 && 
b[28312] == 28312 && 
b[28313] == 28313 && 
b[28314] == 28314 && 
b[28315] == 28315 && 
b[28316] == 28316 && 
b[28317] == 28317 && 
b[28318] == 28318 && 
b[28319] == 28319 && 
b[28320] == 28320 && 
b[28321] == 28321 && 
b[28322] == 28322 && 
b[28323] == 28323 && 
b[28324] == 28324 && 
b[28325] == 28325 && 
b[28326] == 28326 && 
b[28327] == 28327 && 
b[28328] == 28328 && 
b[28329] == 28329 && 
b[28330] == 28330 && 
b[28331] == 28331 && 
b[28332] == 28332 && 
b[28333] == 28333 && 
b[28334] == 28334 && 
b[28335] == 28335 && 
b[28336] == 28336 && 
b[28337] == 28337 && 
b[28338] == 28338 && 
b[28339] == 28339 && 
b[28340] == 28340 && 
b[28341] == 28341 && 
b[28342] == 28342 && 
b[28343] == 28343 && 
b[28344] == 28344 && 
b[28345] == 28345 && 
b[28346] == 28346 && 
b[28347] == 28347 && 
b[28348] == 28348 && 
b[28349] == 28349 && 
b[28350] == 28350 && 
b[28351] == 28351 && 
b[28352] == 28352 && 
b[28353] == 28353 && 
b[28354] == 28354 && 
b[28355] == 28355 && 
b[28356] == 28356 && 
b[28357] == 28357 && 
b[28358] == 28358 && 
b[28359] == 28359 && 
b[28360] == 28360 && 
b[28361] == 28361 && 
b[28362] == 28362 && 
b[28363] == 28363 && 
b[28364] == 28364 && 
b[28365] == 28365 && 
b[28366] == 28366 && 
b[28367] == 28367 && 
b[28368] == 28368 && 
b[28369] == 28369 && 
b[28370] == 28370 && 
b[28371] == 28371 && 
b[28372] == 28372 && 
b[28373] == 28373 && 
b[28374] == 28374 && 
b[28375] == 28375 && 
b[28376] == 28376 && 
b[28377] == 28377 && 
b[28378] == 28378 && 
b[28379] == 28379 && 
b[28380] == 28380 && 
b[28381] == 28381 && 
b[28382] == 28382 && 
b[28383] == 28383 && 
b[28384] == 28384 && 
b[28385] == 28385 && 
b[28386] == 28386 && 
b[28387] == 28387 && 
b[28388] == 28388 && 
b[28389] == 28389 && 
b[28390] == 28390 && 
b[28391] == 28391 && 
b[28392] == 28392 && 
b[28393] == 28393 && 
b[28394] == 28394 && 
b[28395] == 28395 && 
b[28396] == 28396 && 
b[28397] == 28397 && 
b[28398] == 28398 && 
b[28399] == 28399 && 
b[28400] == 28400 && 
b[28401] == 28401 && 
b[28402] == 28402 && 
b[28403] == 28403 && 
b[28404] == 28404 && 
b[28405] == 28405 && 
b[28406] == 28406 && 
b[28407] == 28407 && 
b[28408] == 28408 && 
b[28409] == 28409 && 
b[28410] == 28410 && 
b[28411] == 28411 && 
b[28412] == 28412 && 
b[28413] == 28413 && 
b[28414] == 28414 && 
b[28415] == 28415 && 
b[28416] == 28416 && 
b[28417] == 28417 && 
b[28418] == 28418 && 
b[28419] == 28419 && 
b[28420] == 28420 && 
b[28421] == 28421 && 
b[28422] == 28422 && 
b[28423] == 28423 && 
b[28424] == 28424 && 
b[28425] == 28425 && 
b[28426] == 28426 && 
b[28427] == 28427 && 
b[28428] == 28428 && 
b[28429] == 28429 && 
b[28430] == 28430 && 
b[28431] == 28431 && 
b[28432] == 28432 && 
b[28433] == 28433 && 
b[28434] == 28434 && 
b[28435] == 28435 && 
b[28436] == 28436 && 
b[28437] == 28437 && 
b[28438] == 28438 && 
b[28439] == 28439 && 
b[28440] == 28440 && 
b[28441] == 28441 && 
b[28442] == 28442 && 
b[28443] == 28443 && 
b[28444] == 28444 && 
b[28445] == 28445 && 
b[28446] == 28446 && 
b[28447] == 28447 && 
b[28448] == 28448 && 
b[28449] == 28449 && 
b[28450] == 28450 && 
b[28451] == 28451 && 
b[28452] == 28452 && 
b[28453] == 28453 && 
b[28454] == 28454 && 
b[28455] == 28455 && 
b[28456] == 28456 && 
b[28457] == 28457 && 
b[28458] == 28458 && 
b[28459] == 28459 && 
b[28460] == 28460 && 
b[28461] == 28461 && 
b[28462] == 28462 && 
b[28463] == 28463 && 
b[28464] == 28464 && 
b[28465] == 28465 && 
b[28466] == 28466 && 
b[28467] == 28467 && 
b[28468] == 28468 && 
b[28469] == 28469 && 
b[28470] == 28470 && 
b[28471] == 28471 && 
b[28472] == 28472 && 
b[28473] == 28473 && 
b[28474] == 28474 && 
b[28475] == 28475 && 
b[28476] == 28476 && 
b[28477] == 28477 && 
b[28478] == 28478 && 
b[28479] == 28479 && 
b[28480] == 28480 && 
b[28481] == 28481 && 
b[28482] == 28482 && 
b[28483] == 28483 && 
b[28484] == 28484 && 
b[28485] == 28485 && 
b[28486] == 28486 && 
b[28487] == 28487 && 
b[28488] == 28488 && 
b[28489] == 28489 && 
b[28490] == 28490 && 
b[28491] == 28491 && 
b[28492] == 28492 && 
b[28493] == 28493 && 
b[28494] == 28494 && 
b[28495] == 28495 && 
b[28496] == 28496 && 
b[28497] == 28497 && 
b[28498] == 28498 && 
b[28499] == 28499 && 
b[28500] == 28500 && 
b[28501] == 28501 && 
b[28502] == 28502 && 
b[28503] == 28503 && 
b[28504] == 28504 && 
b[28505] == 28505 && 
b[28506] == 28506 && 
b[28507] == 28507 && 
b[28508] == 28508 && 
b[28509] == 28509 && 
b[28510] == 28510 && 
b[28511] == 28511 && 
b[28512] == 28512 && 
b[28513] == 28513 && 
b[28514] == 28514 && 
b[28515] == 28515 && 
b[28516] == 28516 && 
b[28517] == 28517 && 
b[28518] == 28518 && 
b[28519] == 28519 && 
b[28520] == 28520 && 
b[28521] == 28521 && 
b[28522] == 28522 && 
b[28523] == 28523 && 
b[28524] == 28524 && 
b[28525] == 28525 && 
b[28526] == 28526 && 
b[28527] == 28527 && 
b[28528] == 28528 && 
b[28529] == 28529 && 
b[28530] == 28530 && 
b[28531] == 28531 && 
b[28532] == 28532 && 
b[28533] == 28533 && 
b[28534] == 28534 && 
b[28535] == 28535 && 
b[28536] == 28536 && 
b[28537] == 28537 && 
b[28538] == 28538 && 
b[28539] == 28539 && 
b[28540] == 28540 && 
b[28541] == 28541 && 
b[28542] == 28542 && 
b[28543] == 28543 && 
b[28544] == 28544 && 
b[28545] == 28545 && 
b[28546] == 28546 && 
b[28547] == 28547 && 
b[28548] == 28548 && 
b[28549] == 28549 && 
b[28550] == 28550 && 
b[28551] == 28551 && 
b[28552] == 28552 && 
b[28553] == 28553 && 
b[28554] == 28554 && 
b[28555] == 28555 && 
b[28556] == 28556 && 
b[28557] == 28557 && 
b[28558] == 28558 && 
b[28559] == 28559 && 
b[28560] == 28560 && 
b[28561] == 28561 && 
b[28562] == 28562 && 
b[28563] == 28563 && 
b[28564] == 28564 && 
b[28565] == 28565 && 
b[28566] == 28566 && 
b[28567] == 28567 && 
b[28568] == 28568 && 
b[28569] == 28569 && 
b[28570] == 28570 && 
b[28571] == 28571 && 
b[28572] == 28572 && 
b[28573] == 28573 && 
b[28574] == 28574 && 
b[28575] == 28575 && 
b[28576] == 28576 && 
b[28577] == 28577 && 
b[28578] == 28578 && 
b[28579] == 28579 && 
b[28580] == 28580 && 
b[28581] == 28581 && 
b[28582] == 28582 && 
b[28583] == 28583 && 
b[28584] == 28584 && 
b[28585] == 28585 && 
b[28586] == 28586 && 
b[28587] == 28587 && 
b[28588] == 28588 && 
b[28589] == 28589 && 
b[28590] == 28590 && 
b[28591] == 28591 && 
b[28592] == 28592 && 
b[28593] == 28593 && 
b[28594] == 28594 && 
b[28595] == 28595 && 
b[28596] == 28596 && 
b[28597] == 28597 && 
b[28598] == 28598 && 
b[28599] == 28599 && 
b[28600] == 28600 && 
b[28601] == 28601 && 
b[28602] == 28602 && 
b[28603] == 28603 && 
b[28604] == 28604 && 
b[28605] == 28605 && 
b[28606] == 28606 && 
b[28607] == 28607 && 
b[28608] == 28608 && 
b[28609] == 28609 && 
b[28610] == 28610 && 
b[28611] == 28611 && 
b[28612] == 28612 && 
b[28613] == 28613 && 
b[28614] == 28614 && 
b[28615] == 28615 && 
b[28616] == 28616 && 
b[28617] == 28617 && 
b[28618] == 28618 && 
b[28619] == 28619 && 
b[28620] == 28620 && 
b[28621] == 28621 && 
b[28622] == 28622 && 
b[28623] == 28623 && 
b[28624] == 28624 && 
b[28625] == 28625 && 
b[28626] == 28626 && 
b[28627] == 28627 && 
b[28628] == 28628 && 
b[28629] == 28629 && 
b[28630] == 28630 && 
b[28631] == 28631 && 
b[28632] == 28632 && 
b[28633] == 28633 && 
b[28634] == 28634 && 
b[28635] == 28635 && 
b[28636] == 28636 && 
b[28637] == 28637 && 
b[28638] == 28638 && 
b[28639] == 28639 && 
b[28640] == 28640 && 
b[28641] == 28641 && 
b[28642] == 28642 && 
b[28643] == 28643 && 
b[28644] == 28644 && 
b[28645] == 28645 && 
b[28646] == 28646 && 
b[28647] == 28647 && 
b[28648] == 28648 && 
b[28649] == 28649 && 
b[28650] == 28650 && 
b[28651] == 28651 && 
b[28652] == 28652 && 
b[28653] == 28653 && 
b[28654] == 28654 && 
b[28655] == 28655 && 
b[28656] == 28656 && 
b[28657] == 28657 && 
b[28658] == 28658 && 
b[28659] == 28659 && 
b[28660] == 28660 && 
b[28661] == 28661 && 
b[28662] == 28662 && 
b[28663] == 28663 && 
b[28664] == 28664 && 
b[28665] == 28665 && 
b[28666] == 28666 && 
b[28667] == 28667 && 
b[28668] == 28668 && 
b[28669] == 28669 && 
b[28670] == 28670 && 
b[28671] == 28671 && 
b[28672] == 28672 && 
b[28673] == 28673 && 
b[28674] == 28674 && 
b[28675] == 28675 && 
b[28676] == 28676 && 
b[28677] == 28677 && 
b[28678] == 28678 && 
b[28679] == 28679 && 
b[28680] == 28680 && 
b[28681] == 28681 && 
b[28682] == 28682 && 
b[28683] == 28683 && 
b[28684] == 28684 && 
b[28685] == 28685 && 
b[28686] == 28686 && 
b[28687] == 28687 && 
b[28688] == 28688 && 
b[28689] == 28689 && 
b[28690] == 28690 && 
b[28691] == 28691 && 
b[28692] == 28692 && 
b[28693] == 28693 && 
b[28694] == 28694 && 
b[28695] == 28695 && 
b[28696] == 28696 && 
b[28697] == 28697 && 
b[28698] == 28698 && 
b[28699] == 28699 && 
b[28700] == 28700 && 
b[28701] == 28701 && 
b[28702] == 28702 && 
b[28703] == 28703 && 
b[28704] == 28704 && 
b[28705] == 28705 && 
b[28706] == 28706 && 
b[28707] == 28707 && 
b[28708] == 28708 && 
b[28709] == 28709 && 
b[28710] == 28710 && 
b[28711] == 28711 && 
b[28712] == 28712 && 
b[28713] == 28713 && 
b[28714] == 28714 && 
b[28715] == 28715 && 
b[28716] == 28716 && 
b[28717] == 28717 && 
b[28718] == 28718 && 
b[28719] == 28719 && 
b[28720] == 28720 && 
b[28721] == 28721 && 
b[28722] == 28722 && 
b[28723] == 28723 && 
b[28724] == 28724 && 
b[28725] == 28725 && 
b[28726] == 28726 && 
b[28727] == 28727 && 
b[28728] == 28728 && 
b[28729] == 28729 && 
b[28730] == 28730 && 
b[28731] == 28731 && 
b[28732] == 28732 && 
b[28733] == 28733 && 
b[28734] == 28734 && 
b[28735] == 28735 && 
b[28736] == 28736 && 
b[28737] == 28737 && 
b[28738] == 28738 && 
b[28739] == 28739 && 
b[28740] == 28740 && 
b[28741] == 28741 && 
b[28742] == 28742 && 
b[28743] == 28743 && 
b[28744] == 28744 && 
b[28745] == 28745 && 
b[28746] == 28746 && 
b[28747] == 28747 && 
b[28748] == 28748 && 
b[28749] == 28749 && 
b[28750] == 28750 && 
b[28751] == 28751 && 
b[28752] == 28752 && 
b[28753] == 28753 && 
b[28754] == 28754 && 
b[28755] == 28755 && 
b[28756] == 28756 && 
b[28757] == 28757 && 
b[28758] == 28758 && 
b[28759] == 28759 && 
b[28760] == 28760 && 
b[28761] == 28761 && 
b[28762] == 28762 && 
b[28763] == 28763 && 
b[28764] == 28764 && 
b[28765] == 28765 && 
b[28766] == 28766 && 
b[28767] == 28767 && 
b[28768] == 28768 && 
b[28769] == 28769 && 
b[28770] == 28770 && 
b[28771] == 28771 && 
b[28772] == 28772 && 
b[28773] == 28773 && 
b[28774] == 28774 && 
b[28775] == 28775 && 
b[28776] == 28776 && 
b[28777] == 28777 && 
b[28778] == 28778 && 
b[28779] == 28779 && 
b[28780] == 28780 && 
b[28781] == 28781 && 
b[28782] == 28782 && 
b[28783] == 28783 && 
b[28784] == 28784 && 
b[28785] == 28785 && 
b[28786] == 28786 && 
b[28787] == 28787 && 
b[28788] == 28788 && 
b[28789] == 28789 && 
b[28790] == 28790 && 
b[28791] == 28791 && 
b[28792] == 28792 && 
b[28793] == 28793 && 
b[28794] == 28794 && 
b[28795] == 28795 && 
b[28796] == 28796 && 
b[28797] == 28797 && 
b[28798] == 28798 && 
b[28799] == 28799 && 
b[28800] == 28800 && 
b[28801] == 28801 && 
b[28802] == 28802 && 
b[28803] == 28803 && 
b[28804] == 28804 && 
b[28805] == 28805 && 
b[28806] == 28806 && 
b[28807] == 28807 && 
b[28808] == 28808 && 
b[28809] == 28809 && 
b[28810] == 28810 && 
b[28811] == 28811 && 
b[28812] == 28812 && 
b[28813] == 28813 && 
b[28814] == 28814 && 
b[28815] == 28815 && 
b[28816] == 28816 && 
b[28817] == 28817 && 
b[28818] == 28818 && 
b[28819] == 28819 && 
b[28820] == 28820 && 
b[28821] == 28821 && 
b[28822] == 28822 && 
b[28823] == 28823 && 
b[28824] == 28824 && 
b[28825] == 28825 && 
b[28826] == 28826 && 
b[28827] == 28827 && 
b[28828] == 28828 && 
b[28829] == 28829 && 
b[28830] == 28830 && 
b[28831] == 28831 && 
b[28832] == 28832 && 
b[28833] == 28833 && 
b[28834] == 28834 && 
b[28835] == 28835 && 
b[28836] == 28836 && 
b[28837] == 28837 && 
b[28838] == 28838 && 
b[28839] == 28839 && 
b[28840] == 28840 && 
b[28841] == 28841 && 
b[28842] == 28842 && 
b[28843] == 28843 && 
b[28844] == 28844 && 
b[28845] == 28845 && 
b[28846] == 28846 && 
b[28847] == 28847 && 
b[28848] == 28848 && 
b[28849] == 28849 && 
b[28850] == 28850 && 
b[28851] == 28851 && 
b[28852] == 28852 && 
b[28853] == 28853 && 
b[28854] == 28854 && 
b[28855] == 28855 && 
b[28856] == 28856 && 
b[28857] == 28857 && 
b[28858] == 28858 && 
b[28859] == 28859 && 
b[28860] == 28860 && 
b[28861] == 28861 && 
b[28862] == 28862 && 
b[28863] == 28863 && 
b[28864] == 28864 && 
b[28865] == 28865 && 
b[28866] == 28866 && 
b[28867] == 28867 && 
b[28868] == 28868 && 
b[28869] == 28869 && 
b[28870] == 28870 && 
b[28871] == 28871 && 
b[28872] == 28872 && 
b[28873] == 28873 && 
b[28874] == 28874 && 
b[28875] == 28875 && 
b[28876] == 28876 && 
b[28877] == 28877 && 
b[28878] == 28878 && 
b[28879] == 28879 && 
b[28880] == 28880 && 
b[28881] == 28881 && 
b[28882] == 28882 && 
b[28883] == 28883 && 
b[28884] == 28884 && 
b[28885] == 28885 && 
b[28886] == 28886 && 
b[28887] == 28887 && 
b[28888] == 28888 && 
b[28889] == 28889 && 
b[28890] == 28890 && 
b[28891] == 28891 && 
b[28892] == 28892 && 
b[28893] == 28893 && 
b[28894] == 28894 && 
b[28895] == 28895 && 
b[28896] == 28896 && 
b[28897] == 28897 && 
b[28898] == 28898 && 
b[28899] == 28899 && 
b[28900] == 28900 && 
b[28901] == 28901 && 
b[28902] == 28902 && 
b[28903] == 28903 && 
b[28904] == 28904 && 
b[28905] == 28905 && 
b[28906] == 28906 && 
b[28907] == 28907 && 
b[28908] == 28908 && 
b[28909] == 28909 && 
b[28910] == 28910 && 
b[28911] == 28911 && 
b[28912] == 28912 && 
b[28913] == 28913 && 
b[28914] == 28914 && 
b[28915] == 28915 && 
b[28916] == 28916 && 
b[28917] == 28917 && 
b[28918] == 28918 && 
b[28919] == 28919 && 
b[28920] == 28920 && 
b[28921] == 28921 && 
b[28922] == 28922 && 
b[28923] == 28923 && 
b[28924] == 28924 && 
b[28925] == 28925 && 
b[28926] == 28926 && 
b[28927] == 28927 && 
b[28928] == 28928 && 
b[28929] == 28929 && 
b[28930] == 28930 && 
b[28931] == 28931 && 
b[28932] == 28932 && 
b[28933] == 28933 && 
b[28934] == 28934 && 
b[28935] == 28935 && 
b[28936] == 28936 && 
b[28937] == 28937 && 
b[28938] == 28938 && 
b[28939] == 28939 && 
b[28940] == 28940 && 
b[28941] == 28941 && 
b[28942] == 28942 && 
b[28943] == 28943 && 
b[28944] == 28944 && 
b[28945] == 28945 && 
b[28946] == 28946 && 
b[28947] == 28947 && 
b[28948] == 28948 && 
b[28949] == 28949 && 
b[28950] == 28950 && 
b[28951] == 28951 && 
b[28952] == 28952 && 
b[28953] == 28953 && 
b[28954] == 28954 && 
b[28955] == 28955 && 
b[28956] == 28956 && 
b[28957] == 28957 && 
b[28958] == 28958 && 
b[28959] == 28959 && 
b[28960] == 28960 && 
b[28961] == 28961 && 
b[28962] == 28962 && 
b[28963] == 28963 && 
b[28964] == 28964 && 
b[28965] == 28965 && 
b[28966] == 28966 && 
b[28967] == 28967 && 
b[28968] == 28968 && 
b[28969] == 28969 && 
b[28970] == 28970 && 
b[28971] == 28971 && 
b[28972] == 28972 && 
b[28973] == 28973 && 
b[28974] == 28974 && 
b[28975] == 28975 && 
b[28976] == 28976 && 
b[28977] == 28977 && 
b[28978] == 28978 && 
b[28979] == 28979 && 
b[28980] == 28980 && 
b[28981] == 28981 && 
b[28982] == 28982 && 
b[28983] == 28983 && 
b[28984] == 28984 && 
b[28985] == 28985 && 
b[28986] == 28986 && 
b[28987] == 28987 && 
b[28988] == 28988 && 
b[28989] == 28989 && 
b[28990] == 28990 && 
b[28991] == 28991 && 
b[28992] == 28992 && 
b[28993] == 28993 && 
b[28994] == 28994 && 
b[28995] == 28995 && 
b[28996] == 28996 && 
b[28997] == 28997 && 
b[28998] == 28998 && 
b[28999] == 28999 && 
b[29000] == 29000 && 
b[29001] == 29001 && 
b[29002] == 29002 && 
b[29003] == 29003 && 
b[29004] == 29004 && 
b[29005] == 29005 && 
b[29006] == 29006 && 
b[29007] == 29007 && 
b[29008] == 29008 && 
b[29009] == 29009 && 
b[29010] == 29010 && 
b[29011] == 29011 && 
b[29012] == 29012 && 
b[29013] == 29013 && 
b[29014] == 29014 && 
b[29015] == 29015 && 
b[29016] == 29016 && 
b[29017] == 29017 && 
b[29018] == 29018 && 
b[29019] == 29019 && 
b[29020] == 29020 && 
b[29021] == 29021 && 
b[29022] == 29022 && 
b[29023] == 29023 && 
b[29024] == 29024 && 
b[29025] == 29025 && 
b[29026] == 29026 && 
b[29027] == 29027 && 
b[29028] == 29028 && 
b[29029] == 29029 && 
b[29030] == 29030 && 
b[29031] == 29031 && 
b[29032] == 29032 && 
b[29033] == 29033 && 
b[29034] == 29034 && 
b[29035] == 29035 && 
b[29036] == 29036 && 
b[29037] == 29037 && 
b[29038] == 29038 && 
b[29039] == 29039 && 
b[29040] == 29040 && 
b[29041] == 29041 && 
b[29042] == 29042 && 
b[29043] == 29043 && 
b[29044] == 29044 && 
b[29045] == 29045 && 
b[29046] == 29046 && 
b[29047] == 29047 && 
b[29048] == 29048 && 
b[29049] == 29049 && 
b[29050] == 29050 && 
b[29051] == 29051 && 
b[29052] == 29052 && 
b[29053] == 29053 && 
b[29054] == 29054 && 
b[29055] == 29055 && 
b[29056] == 29056 && 
b[29057] == 29057 && 
b[29058] == 29058 && 
b[29059] == 29059 && 
b[29060] == 29060 && 
b[29061] == 29061 && 
b[29062] == 29062 && 
b[29063] == 29063 && 
b[29064] == 29064 && 
b[29065] == 29065 && 
b[29066] == 29066 && 
b[29067] == 29067 && 
b[29068] == 29068 && 
b[29069] == 29069 && 
b[29070] == 29070 && 
b[29071] == 29071 && 
b[29072] == 29072 && 
b[29073] == 29073 && 
b[29074] == 29074 && 
b[29075] == 29075 && 
b[29076] == 29076 && 
b[29077] == 29077 && 
b[29078] == 29078 && 
b[29079] == 29079 && 
b[29080] == 29080 && 
b[29081] == 29081 && 
b[29082] == 29082 && 
b[29083] == 29083 && 
b[29084] == 29084 && 
b[29085] == 29085 && 
b[29086] == 29086 && 
b[29087] == 29087 && 
b[29088] == 29088 && 
b[29089] == 29089 && 
b[29090] == 29090 && 
b[29091] == 29091 && 
b[29092] == 29092 && 
b[29093] == 29093 && 
b[29094] == 29094 && 
b[29095] == 29095 && 
b[29096] == 29096 && 
b[29097] == 29097 && 
b[29098] == 29098 && 
b[29099] == 29099 && 
b[29100] == 29100 && 
b[29101] == 29101 && 
b[29102] == 29102 && 
b[29103] == 29103 && 
b[29104] == 29104 && 
b[29105] == 29105 && 
b[29106] == 29106 && 
b[29107] == 29107 && 
b[29108] == 29108 && 
b[29109] == 29109 && 
b[29110] == 29110 && 
b[29111] == 29111 && 
b[29112] == 29112 && 
b[29113] == 29113 && 
b[29114] == 29114 && 
b[29115] == 29115 && 
b[29116] == 29116 && 
b[29117] == 29117 && 
b[29118] == 29118 && 
b[29119] == 29119 && 
b[29120] == 29120 && 
b[29121] == 29121 && 
b[29122] == 29122 && 
b[29123] == 29123 && 
b[29124] == 29124 && 
b[29125] == 29125 && 
b[29126] == 29126 && 
b[29127] == 29127 && 
b[29128] == 29128 && 
b[29129] == 29129 && 
b[29130] == 29130 && 
b[29131] == 29131 && 
b[29132] == 29132 && 
b[29133] == 29133 && 
b[29134] == 29134 && 
b[29135] == 29135 && 
b[29136] == 29136 && 
b[29137] == 29137 && 
b[29138] == 29138 && 
b[29139] == 29139 && 
b[29140] == 29140 && 
b[29141] == 29141 && 
b[29142] == 29142 && 
b[29143] == 29143 && 
b[29144] == 29144 && 
b[29145] == 29145 && 
b[29146] == 29146 && 
b[29147] == 29147 && 
b[29148] == 29148 && 
b[29149] == 29149 && 
b[29150] == 29150 && 
b[29151] == 29151 && 
b[29152] == 29152 && 
b[29153] == 29153 && 
b[29154] == 29154 && 
b[29155] == 29155 && 
b[29156] == 29156 && 
b[29157] == 29157 && 
b[29158] == 29158 && 
b[29159] == 29159 && 
b[29160] == 29160 && 
b[29161] == 29161 && 
b[29162] == 29162 && 
b[29163] == 29163 && 
b[29164] == 29164 && 
b[29165] == 29165 && 
b[29166] == 29166 && 
b[29167] == 29167 && 
b[29168] == 29168 && 
b[29169] == 29169 && 
b[29170] == 29170 && 
b[29171] == 29171 && 
b[29172] == 29172 && 
b[29173] == 29173 && 
b[29174] == 29174 && 
b[29175] == 29175 && 
b[29176] == 29176 && 
b[29177] == 29177 && 
b[29178] == 29178 && 
b[29179] == 29179 && 
b[29180] == 29180 && 
b[29181] == 29181 && 
b[29182] == 29182 && 
b[29183] == 29183 && 
b[29184] == 29184 && 
b[29185] == 29185 && 
b[29186] == 29186 && 
b[29187] == 29187 && 
b[29188] == 29188 && 
b[29189] == 29189 && 
b[29190] == 29190 && 
b[29191] == 29191 && 
b[29192] == 29192 && 
b[29193] == 29193 && 
b[29194] == 29194 && 
b[29195] == 29195 && 
b[29196] == 29196 && 
b[29197] == 29197 && 
b[29198] == 29198 && 
b[29199] == 29199 && 
b[29200] == 29200 && 
b[29201] == 29201 && 
b[29202] == 29202 && 
b[29203] == 29203 && 
b[29204] == 29204 && 
b[29205] == 29205 && 
b[29206] == 29206 && 
b[29207] == 29207 && 
b[29208] == 29208 && 
b[29209] == 29209 && 
b[29210] == 29210 && 
b[29211] == 29211 && 
b[29212] == 29212 && 
b[29213] == 29213 && 
b[29214] == 29214 && 
b[29215] == 29215 && 
b[29216] == 29216 && 
b[29217] == 29217 && 
b[29218] == 29218 && 
b[29219] == 29219 && 
b[29220] == 29220 && 
b[29221] == 29221 && 
b[29222] == 29222 && 
b[29223] == 29223 && 
b[29224] == 29224 && 
b[29225] == 29225 && 
b[29226] == 29226 && 
b[29227] == 29227 && 
b[29228] == 29228 && 
b[29229] == 29229 && 
b[29230] == 29230 && 
b[29231] == 29231 && 
b[29232] == 29232 && 
b[29233] == 29233 && 
b[29234] == 29234 && 
b[29235] == 29235 && 
b[29236] == 29236 && 
b[29237] == 29237 && 
b[29238] == 29238 && 
b[29239] == 29239 && 
b[29240] == 29240 && 
b[29241] == 29241 && 
b[29242] == 29242 && 
b[29243] == 29243 && 
b[29244] == 29244 && 
b[29245] == 29245 && 
b[29246] == 29246 && 
b[29247] == 29247 && 
b[29248] == 29248 && 
b[29249] == 29249 && 
b[29250] == 29250 && 
b[29251] == 29251 && 
b[29252] == 29252 && 
b[29253] == 29253 && 
b[29254] == 29254 && 
b[29255] == 29255 && 
b[29256] == 29256 && 
b[29257] == 29257 && 
b[29258] == 29258 && 
b[29259] == 29259 && 
b[29260] == 29260 && 
b[29261] == 29261 && 
b[29262] == 29262 && 
b[29263] == 29263 && 
b[29264] == 29264 && 
b[29265] == 29265 && 
b[29266] == 29266 && 
b[29267] == 29267 && 
b[29268] == 29268 && 
b[29269] == 29269 && 
b[29270] == 29270 && 
b[29271] == 29271 && 
b[29272] == 29272 && 
b[29273] == 29273 && 
b[29274] == 29274 && 
b[29275] == 29275 && 
b[29276] == 29276 && 
b[29277] == 29277 && 
b[29278] == 29278 && 
b[29279] == 29279 && 
b[29280] == 29280 && 
b[29281] == 29281 && 
b[29282] == 29282 && 
b[29283] == 29283 && 
b[29284] == 29284 && 
b[29285] == 29285 && 
b[29286] == 29286 && 
b[29287] == 29287 && 
b[29288] == 29288 && 
b[29289] == 29289 && 
b[29290] == 29290 && 
b[29291] == 29291 && 
b[29292] == 29292 && 
b[29293] == 29293 && 
b[29294] == 29294 && 
b[29295] == 29295 && 
b[29296] == 29296 && 
b[29297] == 29297 && 
b[29298] == 29298 && 
b[29299] == 29299 && 
b[29300] == 29300 && 
b[29301] == 29301 && 
b[29302] == 29302 && 
b[29303] == 29303 && 
b[29304] == 29304 && 
b[29305] == 29305 && 
b[29306] == 29306 && 
b[29307] == 29307 && 
b[29308] == 29308 && 
b[29309] == 29309 && 
b[29310] == 29310 && 
b[29311] == 29311 && 
b[29312] == 29312 && 
b[29313] == 29313 && 
b[29314] == 29314 && 
b[29315] == 29315 && 
b[29316] == 29316 && 
b[29317] == 29317 && 
b[29318] == 29318 && 
b[29319] == 29319 && 
b[29320] == 29320 && 
b[29321] == 29321 && 
b[29322] == 29322 && 
b[29323] == 29323 && 
b[29324] == 29324 && 
b[29325] == 29325 && 
b[29326] == 29326 && 
b[29327] == 29327 && 
b[29328] == 29328 && 
b[29329] == 29329 && 
b[29330] == 29330 && 
b[29331] == 29331 && 
b[29332] == 29332 && 
b[29333] == 29333 && 
b[29334] == 29334 && 
b[29335] == 29335 && 
b[29336] == 29336 && 
b[29337] == 29337 && 
b[29338] == 29338 && 
b[29339] == 29339 && 
b[29340] == 29340 && 
b[29341] == 29341 && 
b[29342] == 29342 && 
b[29343] == 29343 && 
b[29344] == 29344 && 
b[29345] == 29345 && 
b[29346] == 29346 && 
b[29347] == 29347 && 
b[29348] == 29348 && 
b[29349] == 29349 && 
b[29350] == 29350 && 
b[29351] == 29351 && 
b[29352] == 29352 && 
b[29353] == 29353 && 
b[29354] == 29354 && 
b[29355] == 29355 && 
b[29356] == 29356 && 
b[29357] == 29357 && 
b[29358] == 29358 && 
b[29359] == 29359 && 
b[29360] == 29360 && 
b[29361] == 29361 && 
b[29362] == 29362 && 
b[29363] == 29363 && 
b[29364] == 29364 && 
b[29365] == 29365 && 
b[29366] == 29366 && 
b[29367] == 29367 && 
b[29368] == 29368 && 
b[29369] == 29369 && 
b[29370] == 29370 && 
b[29371] == 29371 && 
b[29372] == 29372 && 
b[29373] == 29373 && 
b[29374] == 29374 && 
b[29375] == 29375 && 
b[29376] == 29376 && 
b[29377] == 29377 && 
b[29378] == 29378 && 
b[29379] == 29379 && 
b[29380] == 29380 && 
b[29381] == 29381 && 
b[29382] == 29382 && 
b[29383] == 29383 && 
b[29384] == 29384 && 
b[29385] == 29385 && 
b[29386] == 29386 && 
b[29387] == 29387 && 
b[29388] == 29388 && 
b[29389] == 29389 && 
b[29390] == 29390 && 
b[29391] == 29391 && 
b[29392] == 29392 && 
b[29393] == 29393 && 
b[29394] == 29394 && 
b[29395] == 29395 && 
b[29396] == 29396 && 
b[29397] == 29397 && 
b[29398] == 29398 && 
b[29399] == 29399 && 
b[29400] == 29400 && 
b[29401] == 29401 && 
b[29402] == 29402 && 
b[29403] == 29403 && 
b[29404] == 29404 && 
b[29405] == 29405 && 
b[29406] == 29406 && 
b[29407] == 29407 && 
b[29408] == 29408 && 
b[29409] == 29409 && 
b[29410] == 29410 && 
b[29411] == 29411 && 
b[29412] == 29412 && 
b[29413] == 29413 && 
b[29414] == 29414 && 
b[29415] == 29415 && 
b[29416] == 29416 && 
b[29417] == 29417 && 
b[29418] == 29418 && 
b[29419] == 29419 && 
b[29420] == 29420 && 
b[29421] == 29421 && 
b[29422] == 29422 && 
b[29423] == 29423 && 
b[29424] == 29424 && 
b[29425] == 29425 && 
b[29426] == 29426 && 
b[29427] == 29427 && 
b[29428] == 29428 && 
b[29429] == 29429 && 
b[29430] == 29430 && 
b[29431] == 29431 && 
b[29432] == 29432 && 
b[29433] == 29433 && 
b[29434] == 29434 && 
b[29435] == 29435 && 
b[29436] == 29436 && 
b[29437] == 29437 && 
b[29438] == 29438 && 
b[29439] == 29439 && 
b[29440] == 29440 && 
b[29441] == 29441 && 
b[29442] == 29442 && 
b[29443] == 29443 && 
b[29444] == 29444 && 
b[29445] == 29445 && 
b[29446] == 29446 && 
b[29447] == 29447 && 
b[29448] == 29448 && 
b[29449] == 29449 && 
b[29450] == 29450 && 
b[29451] == 29451 && 
b[29452] == 29452 && 
b[29453] == 29453 && 
b[29454] == 29454 && 
b[29455] == 29455 && 
b[29456] == 29456 && 
b[29457] == 29457 && 
b[29458] == 29458 && 
b[29459] == 29459 && 
b[29460] == 29460 && 
b[29461] == 29461 && 
b[29462] == 29462 && 
b[29463] == 29463 && 
b[29464] == 29464 && 
b[29465] == 29465 && 
b[29466] == 29466 && 
b[29467] == 29467 && 
b[29468] == 29468 && 
b[29469] == 29469 && 
b[29470] == 29470 && 
b[29471] == 29471 && 
b[29472] == 29472 && 
b[29473] == 29473 && 
b[29474] == 29474 && 
b[29475] == 29475 && 
b[29476] == 29476 && 
b[29477] == 29477 && 
b[29478] == 29478 && 
b[29479] == 29479 && 
b[29480] == 29480 && 
b[29481] == 29481 && 
b[29482] == 29482 && 
b[29483] == 29483 && 
b[29484] == 29484 && 
b[29485] == 29485 && 
b[29486] == 29486 && 
b[29487] == 29487 && 
b[29488] == 29488 && 
b[29489] == 29489 && 
b[29490] == 29490 && 
b[29491] == 29491 && 
b[29492] == 29492 && 
b[29493] == 29493 && 
b[29494] == 29494 && 
b[29495] == 29495 && 
b[29496] == 29496 && 
b[29497] == 29497 && 
b[29498] == 29498 && 
b[29499] == 29499 && 
b[29500] == 29500 && 
b[29501] == 29501 && 
b[29502] == 29502 && 
b[29503] == 29503 && 
b[29504] == 29504 && 
b[29505] == 29505 && 
b[29506] == 29506 && 
b[29507] == 29507 && 
b[29508] == 29508 && 
b[29509] == 29509 && 
b[29510] == 29510 && 
b[29511] == 29511 && 
b[29512] == 29512 && 
b[29513] == 29513 && 
b[29514] == 29514 && 
b[29515] == 29515 && 
b[29516] == 29516 && 
b[29517] == 29517 && 
b[29518] == 29518 && 
b[29519] == 29519 && 
b[29520] == 29520 && 
b[29521] == 29521 && 
b[29522] == 29522 && 
b[29523] == 29523 && 
b[29524] == 29524 && 
b[29525] == 29525 && 
b[29526] == 29526 && 
b[29527] == 29527 && 
b[29528] == 29528 && 
b[29529] == 29529 && 
b[29530] == 29530 && 
b[29531] == 29531 && 
b[29532] == 29532 && 
b[29533] == 29533 && 
b[29534] == 29534 && 
b[29535] == 29535 && 
b[29536] == 29536 && 
b[29537] == 29537 && 
b[29538] == 29538 && 
b[29539] == 29539 && 
b[29540] == 29540 && 
b[29541] == 29541 && 
b[29542] == 29542 && 
b[29543] == 29543 && 
b[29544] == 29544 && 
b[29545] == 29545 && 
b[29546] == 29546 && 
b[29547] == 29547 && 
b[29548] == 29548 && 
b[29549] == 29549 && 
b[29550] == 29550 && 
b[29551] == 29551 && 
b[29552] == 29552 && 
b[29553] == 29553 && 
b[29554] == 29554 && 
b[29555] == 29555 && 
b[29556] == 29556 && 
b[29557] == 29557 && 
b[29558] == 29558 && 
b[29559] == 29559 && 
b[29560] == 29560 && 
b[29561] == 29561 && 
b[29562] == 29562 && 
b[29563] == 29563 && 
b[29564] == 29564 && 
b[29565] == 29565 && 
b[29566] == 29566 && 
b[29567] == 29567 && 
b[29568] == 29568 && 
b[29569] == 29569 && 
b[29570] == 29570 && 
b[29571] == 29571 && 
b[29572] == 29572 && 
b[29573] == 29573 && 
b[29574] == 29574 && 
b[29575] == 29575 && 
b[29576] == 29576 && 
b[29577] == 29577 && 
b[29578] == 29578 && 
b[29579] == 29579 && 
b[29580] == 29580 && 
b[29581] == 29581 && 
b[29582] == 29582 && 
b[29583] == 29583 && 
b[29584] == 29584 && 
b[29585] == 29585 && 
b[29586] == 29586 && 
b[29587] == 29587 && 
b[29588] == 29588 && 
b[29589] == 29589 && 
b[29590] == 29590 && 
b[29591] == 29591 && 
b[29592] == 29592 && 
b[29593] == 29593 && 
b[29594] == 29594 && 
b[29595] == 29595 && 
b[29596] == 29596 && 
b[29597] == 29597 && 
b[29598] == 29598 && 
b[29599] == 29599 && 
b[29600] == 29600 && 
b[29601] == 29601 && 
b[29602] == 29602 && 
b[29603] == 29603 && 
b[29604] == 29604 && 
b[29605] == 29605 && 
b[29606] == 29606 && 
b[29607] == 29607 && 
b[29608] == 29608 && 
b[29609] == 29609 && 
b[29610] == 29610 && 
b[29611] == 29611 && 
b[29612] == 29612 && 
b[29613] == 29613 && 
b[29614] == 29614 && 
b[29615] == 29615 && 
b[29616] == 29616 && 
b[29617] == 29617 && 
b[29618] == 29618 && 
b[29619] == 29619 && 
b[29620] == 29620 && 
b[29621] == 29621 && 
b[29622] == 29622 && 
b[29623] == 29623 && 
b[29624] == 29624 && 
b[29625] == 29625 && 
b[29626] == 29626 && 
b[29627] == 29627 && 
b[29628] == 29628 && 
b[29629] == 29629 && 
b[29630] == 29630 && 
b[29631] == 29631 && 
b[29632] == 29632 && 
b[29633] == 29633 && 
b[29634] == 29634 && 
b[29635] == 29635 && 
b[29636] == 29636 && 
b[29637] == 29637 && 
b[29638] == 29638 && 
b[29639] == 29639 && 
b[29640] == 29640 && 
b[29641] == 29641 && 
b[29642] == 29642 && 
b[29643] == 29643 && 
b[29644] == 29644 && 
b[29645] == 29645 && 
b[29646] == 29646 && 
b[29647] == 29647 && 
b[29648] == 29648 && 
b[29649] == 29649 && 
b[29650] == 29650 && 
b[29651] == 29651 && 
b[29652] == 29652 && 
b[29653] == 29653 && 
b[29654] == 29654 && 
b[29655] == 29655 && 
b[29656] == 29656 && 
b[29657] == 29657 && 
b[29658] == 29658 && 
b[29659] == 29659 && 
b[29660] == 29660 && 
b[29661] == 29661 && 
b[29662] == 29662 && 
b[29663] == 29663 && 
b[29664] == 29664 && 
b[29665] == 29665 && 
b[29666] == 29666 && 
b[29667] == 29667 && 
b[29668] == 29668 && 
b[29669] == 29669 && 
b[29670] == 29670 && 
b[29671] == 29671 && 
b[29672] == 29672 && 
b[29673] == 29673 && 
b[29674] == 29674 && 
b[29675] == 29675 && 
b[29676] == 29676 && 
b[29677] == 29677 && 
b[29678] == 29678 && 
b[29679] == 29679 && 
b[29680] == 29680 && 
b[29681] == 29681 && 
b[29682] == 29682 && 
b[29683] == 29683 && 
b[29684] == 29684 && 
b[29685] == 29685 && 
b[29686] == 29686 && 
b[29687] == 29687 && 
b[29688] == 29688 && 
b[29689] == 29689 && 
b[29690] == 29690 && 
b[29691] == 29691 && 
b[29692] == 29692 && 
b[29693] == 29693 && 
b[29694] == 29694 && 
b[29695] == 29695 && 
b[29696] == 29696 && 
b[29697] == 29697 && 
b[29698] == 29698 && 
b[29699] == 29699 && 
b[29700] == 29700 && 
b[29701] == 29701 && 
b[29702] == 29702 && 
b[29703] == 29703 && 
b[29704] == 29704 && 
b[29705] == 29705 && 
b[29706] == 29706 && 
b[29707] == 29707 && 
b[29708] == 29708 && 
b[29709] == 29709 && 
b[29710] == 29710 && 
b[29711] == 29711 && 
b[29712] == 29712 && 
b[29713] == 29713 && 
b[29714] == 29714 && 
b[29715] == 29715 && 
b[29716] == 29716 && 
b[29717] == 29717 && 
b[29718] == 29718 && 
b[29719] == 29719 && 
b[29720] == 29720 && 
b[29721] == 29721 && 
b[29722] == 29722 && 
b[29723] == 29723 && 
b[29724] == 29724 && 
b[29725] == 29725 && 
b[29726] == 29726 && 
b[29727] == 29727 && 
b[29728] == 29728 && 
b[29729] == 29729 && 
b[29730] == 29730 && 
b[29731] == 29731 && 
b[29732] == 29732 && 
b[29733] == 29733 && 
b[29734] == 29734 && 
b[29735] == 29735 && 
b[29736] == 29736 && 
b[29737] == 29737 && 
b[29738] == 29738 && 
b[29739] == 29739 && 
b[29740] == 29740 && 
b[29741] == 29741 && 
b[29742] == 29742 && 
b[29743] == 29743 && 
b[29744] == 29744 && 
b[29745] == 29745 && 
b[29746] == 29746 && 
b[29747] == 29747 && 
b[29748] == 29748 && 
b[29749] == 29749 && 
b[29750] == 29750 && 
b[29751] == 29751 && 
b[29752] == 29752 && 
b[29753] == 29753 && 
b[29754] == 29754 && 
b[29755] == 29755 && 
b[29756] == 29756 && 
b[29757] == 29757 && 
b[29758] == 29758 && 
b[29759] == 29759 && 
b[29760] == 29760 && 
b[29761] == 29761 && 
b[29762] == 29762 && 
b[29763] == 29763 && 
b[29764] == 29764 && 
b[29765] == 29765 && 
b[29766] == 29766 && 
b[29767] == 29767 && 
b[29768] == 29768 && 
b[29769] == 29769 && 
b[29770] == 29770 && 
b[29771] == 29771 && 
b[29772] == 29772 && 
b[29773] == 29773 && 
b[29774] == 29774 && 
b[29775] == 29775 && 
b[29776] == 29776 && 
b[29777] == 29777 && 
b[29778] == 29778 && 
b[29779] == 29779 && 
b[29780] == 29780 && 
b[29781] == 29781 && 
b[29782] == 29782 && 
b[29783] == 29783 && 
b[29784] == 29784 && 
b[29785] == 29785 && 
b[29786] == 29786 && 
b[29787] == 29787 && 
b[29788] == 29788 && 
b[29789] == 29789 && 
b[29790] == 29790 && 
b[29791] == 29791 && 
b[29792] == 29792 && 
b[29793] == 29793 && 
b[29794] == 29794 && 
b[29795] == 29795 && 
b[29796] == 29796 && 
b[29797] == 29797 && 
b[29798] == 29798 && 
b[29799] == 29799 && 
b[29800] == 29800 && 
b[29801] == 29801 && 
b[29802] == 29802 && 
b[29803] == 29803 && 
b[29804] == 29804 && 
b[29805] == 29805 && 
b[29806] == 29806 && 
b[29807] == 29807 && 
b[29808] == 29808 && 
b[29809] == 29809 && 
b[29810] == 29810 && 
b[29811] == 29811 && 
b[29812] == 29812 && 
b[29813] == 29813 && 
b[29814] == 29814 && 
b[29815] == 29815 && 
b[29816] == 29816 && 
b[29817] == 29817 && 
b[29818] == 29818 && 
b[29819] == 29819 && 
b[29820] == 29820 && 
b[29821] == 29821 && 
b[29822] == 29822 && 
b[29823] == 29823 && 
b[29824] == 29824 && 
b[29825] == 29825 && 
b[29826] == 29826 && 
b[29827] == 29827 && 
b[29828] == 29828 && 
b[29829] == 29829 && 
b[29830] == 29830 && 
b[29831] == 29831 && 
b[29832] == 29832 && 
b[29833] == 29833 && 
b[29834] == 29834 && 
b[29835] == 29835 && 
b[29836] == 29836 && 
b[29837] == 29837 && 
b[29838] == 29838 && 
b[29839] == 29839 && 
b[29840] == 29840 && 
b[29841] == 29841 && 
b[29842] == 29842 && 
b[29843] == 29843 && 
b[29844] == 29844 && 
b[29845] == 29845 && 
b[29846] == 29846 && 
b[29847] == 29847 && 
b[29848] == 29848 && 
b[29849] == 29849 && 
b[29850] == 29850 && 
b[29851] == 29851 && 
b[29852] == 29852 && 
b[29853] == 29853 && 
b[29854] == 29854 && 
b[29855] == 29855 && 
b[29856] == 29856 && 
b[29857] == 29857 && 
b[29858] == 29858 && 
b[29859] == 29859 && 
b[29860] == 29860 && 
b[29861] == 29861 && 
b[29862] == 29862 && 
b[29863] == 29863 && 
b[29864] == 29864 && 
b[29865] == 29865 && 
b[29866] == 29866 && 
b[29867] == 29867 && 
b[29868] == 29868 && 
b[29869] == 29869 && 
b[29870] == 29870 && 
b[29871] == 29871 && 
b[29872] == 29872 && 
b[29873] == 29873 && 
b[29874] == 29874 && 
b[29875] == 29875 && 
b[29876] == 29876 && 
b[29877] == 29877 && 
b[29878] == 29878 && 
b[29879] == 29879 && 
b[29880] == 29880 && 
b[29881] == 29881 && 
b[29882] == 29882 && 
b[29883] == 29883 && 
b[29884] == 29884 && 
b[29885] == 29885 && 
b[29886] == 29886 && 
b[29887] == 29887 && 
b[29888] == 29888 && 
b[29889] == 29889 && 
b[29890] == 29890 && 
b[29891] == 29891 && 
b[29892] == 29892 && 
b[29893] == 29893 && 
b[29894] == 29894 && 
b[29895] == 29895 && 
b[29896] == 29896 && 
b[29897] == 29897 && 
b[29898] == 29898 && 
b[29899] == 29899 && 
b[29900] == 29900 && 
b[29901] == 29901 && 
b[29902] == 29902 && 
b[29903] == 29903 && 
b[29904] == 29904 && 
b[29905] == 29905 && 
b[29906] == 29906 && 
b[29907] == 29907 && 
b[29908] == 29908 && 
b[29909] == 29909 && 
b[29910] == 29910 && 
b[29911] == 29911 && 
b[29912] == 29912 && 
b[29913] == 29913 && 
b[29914] == 29914 && 
b[29915] == 29915 && 
b[29916] == 29916 && 
b[29917] == 29917 && 
b[29918] == 29918 && 
b[29919] == 29919 && 
b[29920] == 29920 && 
b[29921] == 29921 && 
b[29922] == 29922 && 
b[29923] == 29923 && 
b[29924] == 29924 && 
b[29925] == 29925 && 
b[29926] == 29926 && 
b[29927] == 29927 && 
b[29928] == 29928 && 
b[29929] == 29929 && 
b[29930] == 29930 && 
b[29931] == 29931 && 
b[29932] == 29932 && 
b[29933] == 29933 && 
b[29934] == 29934 && 
b[29935] == 29935 && 
b[29936] == 29936 && 
b[29937] == 29937 && 
b[29938] == 29938 && 
b[29939] == 29939 && 
b[29940] == 29940 && 
b[29941] == 29941 && 
b[29942] == 29942 && 
b[29943] == 29943 && 
b[29944] == 29944 && 
b[29945] == 29945 && 
b[29946] == 29946 && 
b[29947] == 29947 && 
b[29948] == 29948 && 
b[29949] == 29949 && 
b[29950] == 29950 && 
b[29951] == 29951 && 
b[29952] == 29952 && 
b[29953] == 29953 && 
b[29954] == 29954 && 
b[29955] == 29955 && 
b[29956] == 29956 && 
b[29957] == 29957 && 
b[29958] == 29958 && 
b[29959] == 29959 && 
b[29960] == 29960 && 
b[29961] == 29961 && 
b[29962] == 29962 && 
b[29963] == 29963 && 
b[29964] == 29964 && 
b[29965] == 29965 && 
b[29966] == 29966 && 
b[29967] == 29967 && 
b[29968] == 29968 && 
b[29969] == 29969 && 
b[29970] == 29970 && 
b[29971] == 29971 && 
b[29972] == 29972 && 
b[29973] == 29973 && 
b[29974] == 29974 && 
b[29975] == 29975 && 
b[29976] == 29976 && 
b[29977] == 29977 && 
b[29978] == 29978 && 
b[29979] == 29979 && 
b[29980] == 29980 && 
b[29981] == 29981 && 
b[29982] == 29982 && 
b[29983] == 29983 && 
b[29984] == 29984 && 
b[29985] == 29985 && 
b[29986] == 29986 && 
b[29987] == 29987 && 
b[29988] == 29988 && 
b[29989] == 29989 && 
b[29990] == 29990 && 
b[29991] == 29991 && 
b[29992] == 29992 && 
b[29993] == 29993 && 
b[29994] == 29994 && 
b[29995] == 29995 && 
b[29996] == 29996 && 
b[29997] == 29997 && 
b[29998] == 29998 && 
b[29999] == 29999 && 
b[30000] == 30000 && 
b[30001] == 30001 && 
b[30002] == 30002 && 
b[30003] == 30003 && 
b[30004] == 30004 && 
b[30005] == 30005 && 
b[30006] == 30006 && 
b[30007] == 30007 && 
b[30008] == 30008 && 
b[30009] == 30009 && 
b[30010] == 30010 && 
b[30011] == 30011 && 
b[30012] == 30012 && 
b[30013] == 30013 && 
b[30014] == 30014 && 
b[30015] == 30015 && 
b[30016] == 30016 && 
b[30017] == 30017 && 
b[30018] == 30018 && 
b[30019] == 30019 && 
b[30020] == 30020 && 
b[30021] == 30021 && 
b[30022] == 30022 && 
b[30023] == 30023 && 
b[30024] == 30024 && 
b[30025] == 30025 && 
b[30026] == 30026 && 
b[30027] == 30027 && 
b[30028] == 30028 && 
b[30029] == 30029 && 
b[30030] == 30030 && 
b[30031] == 30031 && 
b[30032] == 30032 && 
b[30033] == 30033 && 
b[30034] == 30034 && 
b[30035] == 30035 && 
b[30036] == 30036 && 
b[30037] == 30037 && 
b[30038] == 30038 && 
b[30039] == 30039 && 
b[30040] == 30040 && 
b[30041] == 30041 && 
b[30042] == 30042 && 
b[30043] == 30043 && 
b[30044] == 30044 && 
b[30045] == 30045 && 
b[30046] == 30046 && 
b[30047] == 30047 && 
b[30048] == 30048 && 
b[30049] == 30049 && 
b[30050] == 30050 && 
b[30051] == 30051 && 
b[30052] == 30052 && 
b[30053] == 30053 && 
b[30054] == 30054 && 
b[30055] == 30055 && 
b[30056] == 30056 && 
b[30057] == 30057 && 
b[30058] == 30058 && 
b[30059] == 30059 && 
b[30060] == 30060 && 
b[30061] == 30061 && 
b[30062] == 30062 && 
b[30063] == 30063 && 
b[30064] == 30064 && 
b[30065] == 30065 && 
b[30066] == 30066 && 
b[30067] == 30067 && 
b[30068] == 30068 && 
b[30069] == 30069 && 
b[30070] == 30070 && 
b[30071] == 30071 && 
b[30072] == 30072 && 
b[30073] == 30073 && 
b[30074] == 30074 && 
b[30075] == 30075 && 
b[30076] == 30076 && 
b[30077] == 30077 && 
b[30078] == 30078 && 
b[30079] == 30079 && 
b[30080] == 30080 && 
b[30081] == 30081 && 
b[30082] == 30082 && 
b[30083] == 30083 && 
b[30084] == 30084 && 
b[30085] == 30085 && 
b[30086] == 30086 && 
b[30087] == 30087 && 
b[30088] == 30088 && 
b[30089] == 30089 && 
b[30090] == 30090 && 
b[30091] == 30091 && 
b[30092] == 30092 && 
b[30093] == 30093 && 
b[30094] == 30094 && 
b[30095] == 30095 && 
b[30096] == 30096 && 
b[30097] == 30097 && 
b[30098] == 30098 && 
b[30099] == 30099 && 
b[30100] == 30100 && 
b[30101] == 30101 && 
b[30102] == 30102 && 
b[30103] == 30103 && 
b[30104] == 30104 && 
b[30105] == 30105 && 
b[30106] == 30106 && 
b[30107] == 30107 && 
b[30108] == 30108 && 
b[30109] == 30109 && 
b[30110] == 30110 && 
b[30111] == 30111 && 
b[30112] == 30112 && 
b[30113] == 30113 && 
b[30114] == 30114 && 
b[30115] == 30115 && 
b[30116] == 30116 && 
b[30117] == 30117 && 
b[30118] == 30118 && 
b[30119] == 30119 && 
b[30120] == 30120 && 
b[30121] == 30121 && 
b[30122] == 30122 && 
b[30123] == 30123 && 
b[30124] == 30124 && 
b[30125] == 30125 && 
b[30126] == 30126 && 
b[30127] == 30127 && 
b[30128] == 30128 && 
b[30129] == 30129 && 
b[30130] == 30130 && 
b[30131] == 30131 && 
b[30132] == 30132 && 
b[30133] == 30133 && 
b[30134] == 30134 && 
b[30135] == 30135 && 
b[30136] == 30136 && 
b[30137] == 30137 && 
b[30138] == 30138 && 
b[30139] == 30139 && 
b[30140] == 30140 && 
b[30141] == 30141 && 
b[30142] == 30142 && 
b[30143] == 30143 && 
b[30144] == 30144 && 
b[30145] == 30145 && 
b[30146] == 30146 && 
b[30147] == 30147 && 
b[30148] == 30148 && 
b[30149] == 30149 && 
b[30150] == 30150 && 
b[30151] == 30151 && 
b[30152] == 30152 && 
b[30153] == 30153 && 
b[30154] == 30154 && 
b[30155] == 30155 && 
b[30156] == 30156 && 
b[30157] == 30157 && 
b[30158] == 30158 && 
b[30159] == 30159 && 
b[30160] == 30160 && 
b[30161] == 30161 && 
b[30162] == 30162 && 
b[30163] == 30163 && 
b[30164] == 30164 && 
b[30165] == 30165 && 
b[30166] == 30166 && 
b[30167] == 30167 && 
b[30168] == 30168 && 
b[30169] == 30169 && 
b[30170] == 30170 && 
b[30171] == 30171 && 
b[30172] == 30172 && 
b[30173] == 30173 && 
b[30174] == 30174 && 
b[30175] == 30175 && 
b[30176] == 30176 && 
b[30177] == 30177 && 
b[30178] == 30178 && 
b[30179] == 30179 && 
b[30180] == 30180 && 
b[30181] == 30181 && 
b[30182] == 30182 && 
b[30183] == 30183 && 
b[30184] == 30184 && 
b[30185] == 30185 && 
b[30186] == 30186 && 
b[30187] == 30187 && 
b[30188] == 30188 && 
b[30189] == 30189 && 
b[30190] == 30190 && 
b[30191] == 30191 && 
b[30192] == 30192 && 
b[30193] == 30193 && 
b[30194] == 30194 && 
b[30195] == 30195 && 
b[30196] == 30196 && 
b[30197] == 30197 && 
b[30198] == 30198 && 
b[30199] == 30199 && 
b[30200] == 30200 && 
b[30201] == 30201 && 
b[30202] == 30202 && 
b[30203] == 30203 && 
b[30204] == 30204 && 
b[30205] == 30205 && 
b[30206] == 30206 && 
b[30207] == 30207 && 
b[30208] == 30208 && 
b[30209] == 30209 && 
b[30210] == 30210 && 
b[30211] == 30211 && 
b[30212] == 30212 && 
b[30213] == 30213 && 
b[30214] == 30214 && 
b[30215] == 30215 && 
b[30216] == 30216 && 
b[30217] == 30217 && 
b[30218] == 30218 && 
b[30219] == 30219 && 
b[30220] == 30220 && 
b[30221] == 30221 && 
b[30222] == 30222 && 
b[30223] == 30223 && 
b[30224] == 30224 && 
b[30225] == 30225 && 
b[30226] == 30226 && 
b[30227] == 30227 && 
b[30228] == 30228 && 
b[30229] == 30229 && 
b[30230] == 30230 && 
b[30231] == 30231 && 
b[30232] == 30232 && 
b[30233] == 30233 && 
b[30234] == 30234 && 
b[30235] == 30235 && 
b[30236] == 30236 && 
b[30237] == 30237 && 
b[30238] == 30238 && 
b[30239] == 30239 && 
b[30240] == 30240 && 
b[30241] == 30241 && 
b[30242] == 30242 && 
b[30243] == 30243 && 
b[30244] == 30244 && 
b[30245] == 30245 && 
b[30246] == 30246 && 
b[30247] == 30247 && 
b[30248] == 30248 && 
b[30249] == 30249 && 
b[30250] == 30250 && 
b[30251] == 30251 && 
b[30252] == 30252 && 
b[30253] == 30253 && 
b[30254] == 30254 && 
b[30255] == 30255 && 
b[30256] == 30256 && 
b[30257] == 30257 && 
b[30258] == 30258 && 
b[30259] == 30259 && 
b[30260] == 30260 && 
b[30261] == 30261 && 
b[30262] == 30262 && 
b[30263] == 30263 && 
b[30264] == 30264 && 
b[30265] == 30265 && 
b[30266] == 30266 && 
b[30267] == 30267 && 
b[30268] == 30268 && 
b[30269] == 30269 && 
b[30270] == 30270 && 
b[30271] == 30271 && 
b[30272] == 30272 && 
b[30273] == 30273 && 
b[30274] == 30274 && 
b[30275] == 30275 && 
b[30276] == 30276 && 
b[30277] == 30277 && 
b[30278] == 30278 && 
b[30279] == 30279 && 
b[30280] == 30280 && 
b[30281] == 30281 && 
b[30282] == 30282 && 
b[30283] == 30283 && 
b[30284] == 30284 && 
b[30285] == 30285 && 
b[30286] == 30286 && 
b[30287] == 30287 && 
b[30288] == 30288 && 
b[30289] == 30289 && 
b[30290] == 30290 && 
b[30291] == 30291 && 
b[30292] == 30292 && 
b[30293] == 30293 && 
b[30294] == 30294 && 
b[30295] == 30295 && 
b[30296] == 30296 && 
b[30297] == 30297 && 
b[30298] == 30298 && 
b[30299] == 30299 && 
b[30300] == 30300 && 
b[30301] == 30301 && 
b[30302] == 30302 && 
b[30303] == 30303 && 
b[30304] == 30304 && 
b[30305] == 30305 && 
b[30306] == 30306 && 
b[30307] == 30307 && 
b[30308] == 30308 && 
b[30309] == 30309 && 
b[30310] == 30310 && 
b[30311] == 30311 && 
b[30312] == 30312 && 
b[30313] == 30313 && 
b[30314] == 30314 && 
b[30315] == 30315 && 
b[30316] == 30316 && 
b[30317] == 30317 && 
b[30318] == 30318 && 
b[30319] == 30319 && 
b[30320] == 30320 && 
b[30321] == 30321 && 
b[30322] == 30322 && 
b[30323] == 30323 && 
b[30324] == 30324 && 
b[30325] == 30325 && 
b[30326] == 30326 && 
b[30327] == 30327 && 
b[30328] == 30328 && 
b[30329] == 30329 && 
b[30330] == 30330 && 
b[30331] == 30331 && 
b[30332] == 30332 && 
b[30333] == 30333 && 
b[30334] == 30334 && 
b[30335] == 30335 && 
b[30336] == 30336 && 
b[30337] == 30337 && 
b[30338] == 30338 && 
b[30339] == 30339 && 
b[30340] == 30340 && 
b[30341] == 30341 && 
b[30342] == 30342 && 
b[30343] == 30343 && 
b[30344] == 30344 && 
b[30345] == 30345 && 
b[30346] == 30346 && 
b[30347] == 30347 && 
b[30348] == 30348 && 
b[30349] == 30349 && 
b[30350] == 30350 && 
b[30351] == 30351 && 
b[30352] == 30352 && 
b[30353] == 30353 && 
b[30354] == 30354 && 
b[30355] == 30355 && 
b[30356] == 30356 && 
b[30357] == 30357 && 
b[30358] == 30358 && 
b[30359] == 30359 && 
b[30360] == 30360 && 
b[30361] == 30361 && 
b[30362] == 30362 && 
b[30363] == 30363 && 
b[30364] == 30364 && 
b[30365] == 30365 && 
b[30366] == 30366 && 
b[30367] == 30367 && 
b[30368] == 30368 && 
b[30369] == 30369 && 
b[30370] == 30370 && 
b[30371] == 30371 && 
b[30372] == 30372 && 
b[30373] == 30373 && 
b[30374] == 30374 && 
b[30375] == 30375 && 
b[30376] == 30376 && 
b[30377] == 30377 && 
b[30378] == 30378 && 
b[30379] == 30379 && 
b[30380] == 30380 && 
b[30381] == 30381 && 
b[30382] == 30382 && 
b[30383] == 30383 && 
b[30384] == 30384 && 
b[30385] == 30385 && 
b[30386] == 30386 && 
b[30387] == 30387 && 
b[30388] == 30388 && 
b[30389] == 30389 && 
b[30390] == 30390 && 
b[30391] == 30391 && 
b[30392] == 30392 && 
b[30393] == 30393 && 
b[30394] == 30394 && 
b[30395] == 30395 && 
b[30396] == 30396 && 
b[30397] == 30397 && 
b[30398] == 30398 && 
b[30399] == 30399 && 
b[30400] == 30400 && 
b[30401] == 30401 && 
b[30402] == 30402 && 
b[30403] == 30403 && 
b[30404] == 30404 && 
b[30405] == 30405 && 
b[30406] == 30406 && 
b[30407] == 30407 && 
b[30408] == 30408 && 
b[30409] == 30409 && 
b[30410] == 30410 && 
b[30411] == 30411 && 
b[30412] == 30412 && 
b[30413] == 30413 && 
b[30414] == 30414 && 
b[30415] == 30415 && 
b[30416] == 30416 && 
b[30417] == 30417 && 
b[30418] == 30418 && 
b[30419] == 30419 && 
b[30420] == 30420 && 
b[30421] == 30421 && 
b[30422] == 30422 && 
b[30423] == 30423 && 
b[30424] == 30424 && 
b[30425] == 30425 && 
b[30426] == 30426 && 
b[30427] == 30427 && 
b[30428] == 30428 && 
b[30429] == 30429 && 
b[30430] == 30430 && 
b[30431] == 30431 && 
b[30432] == 30432 && 
b[30433] == 30433 && 
b[30434] == 30434 && 
b[30435] == 30435 && 
b[30436] == 30436 && 
b[30437] == 30437 && 
b[30438] == 30438 && 
b[30439] == 30439 && 
b[30440] == 30440 && 
b[30441] == 30441 && 
b[30442] == 30442 && 
b[30443] == 30443 && 
b[30444] == 30444 && 
b[30445] == 30445 && 
b[30446] == 30446 && 
b[30447] == 30447 && 
b[30448] == 30448 && 
b[30449] == 30449 && 
b[30450] == 30450 && 
b[30451] == 30451 && 
b[30452] == 30452 && 
b[30453] == 30453 && 
b[30454] == 30454 && 
b[30455] == 30455 && 
b[30456] == 30456 && 
b[30457] == 30457 && 
b[30458] == 30458 && 
b[30459] == 30459 && 
b[30460] == 30460 && 
b[30461] == 30461 && 
b[30462] == 30462 && 
b[30463] == 30463 && 
b[30464] == 30464 && 
b[30465] == 30465 && 
b[30466] == 30466 && 
b[30467] == 30467 && 
b[30468] == 30468 && 
b[30469] == 30469 && 
b[30470] == 30470 && 
b[30471] == 30471 && 
b[30472] == 30472 && 
b[30473] == 30473 && 
b[30474] == 30474 && 
b[30475] == 30475 && 
b[30476] == 30476 && 
b[30477] == 30477 && 
b[30478] == 30478 && 
b[30479] == 30479 && 
b[30480] == 30480 && 
b[30481] == 30481 && 
b[30482] == 30482 && 
b[30483] == 30483 && 
b[30484] == 30484 && 
b[30485] == 30485 && 
b[30486] == 30486 && 
b[30487] == 30487 && 
b[30488] == 30488 && 
b[30489] == 30489 && 
b[30490] == 30490 && 
b[30491] == 30491 && 
b[30492] == 30492 && 
b[30493] == 30493 && 
b[30494] == 30494 && 
b[30495] == 30495 && 
b[30496] == 30496 && 
b[30497] == 30497 && 
b[30498] == 30498 && 
b[30499] == 30499 && 
b[30500] == 30500 && 
b[30501] == 30501 && 
b[30502] == 30502 && 
b[30503] == 30503 && 
b[30504] == 30504 && 
b[30505] == 30505 && 
b[30506] == 30506 && 
b[30507] == 30507 && 
b[30508] == 30508 && 
b[30509] == 30509 && 
b[30510] == 30510 && 
b[30511] == 30511 && 
b[30512] == 30512 && 
b[30513] == 30513 && 
b[30514] == 30514 && 
b[30515] == 30515 && 
b[30516] == 30516 && 
b[30517] == 30517 && 
b[30518] == 30518 && 
b[30519] == 30519 && 
b[30520] == 30520 && 
b[30521] == 30521 && 
b[30522] == 30522 && 
b[30523] == 30523 && 
b[30524] == 30524 && 
b[30525] == 30525 && 
b[30526] == 30526 && 
b[30527] == 30527 && 
b[30528] == 30528 && 
b[30529] == 30529 && 
b[30530] == 30530 && 
b[30531] == 30531 && 
b[30532] == 30532 && 
b[30533] == 30533 && 
b[30534] == 30534 && 
b[30535] == 30535 && 
b[30536] == 30536 && 
b[30537] == 30537 && 
b[30538] == 30538 && 
b[30539] == 30539 && 
b[30540] == 30540 && 
b[30541] == 30541 && 
b[30542] == 30542 && 
b[30543] == 30543 && 
b[30544] == 30544 && 
b[30545] == 30545 && 
b[30546] == 30546 && 
b[30547] == 30547 && 
b[30548] == 30548 && 
b[30549] == 30549 && 
b[30550] == 30550 && 
b[30551] == 30551 && 
b[30552] == 30552 && 
b[30553] == 30553 && 
b[30554] == 30554 && 
b[30555] == 30555 && 
b[30556] == 30556 && 
b[30557] == 30557 && 
b[30558] == 30558 && 
b[30559] == 30559 && 
b[30560] == 30560 && 
b[30561] == 30561 && 
b[30562] == 30562 && 
b[30563] == 30563 && 
b[30564] == 30564 && 
b[30565] == 30565 && 
b[30566] == 30566 && 
b[30567] == 30567 && 
b[30568] == 30568 && 
b[30569] == 30569 && 
b[30570] == 30570 && 
b[30571] == 30571 && 
b[30572] == 30572 && 
b[30573] == 30573 && 
b[30574] == 30574 && 
b[30575] == 30575 && 
b[30576] == 30576 && 
b[30577] == 30577 && 
b[30578] == 30578 && 
b[30579] == 30579 && 
b[30580] == 30580 && 
b[30581] == 30581 && 
b[30582] == 30582 && 
b[30583] == 30583 && 
b[30584] == 30584 && 
b[30585] == 30585 && 
b[30586] == 30586 && 
b[30587] == 30587 && 
b[30588] == 30588 && 
b[30589] == 30589 && 
b[30590] == 30590 && 
b[30591] == 30591 && 
b[30592] == 30592 && 
b[30593] == 30593 && 
b[30594] == 30594 && 
b[30595] == 30595 && 
b[30596] == 30596 && 
b[30597] == 30597 && 
b[30598] == 30598 && 
b[30599] == 30599 && 
b[30600] == 30600 && 
b[30601] == 30601 && 
b[30602] == 30602 && 
b[30603] == 30603 && 
b[30604] == 30604 && 
b[30605] == 30605 && 
b[30606] == 30606 && 
b[30607] == 30607 && 
b[30608] == 30608 && 
b[30609] == 30609 && 
b[30610] == 30610 && 
b[30611] == 30611 && 
b[30612] == 30612 && 
b[30613] == 30613 && 
b[30614] == 30614 && 
b[30615] == 30615 && 
b[30616] == 30616 && 
b[30617] == 30617 && 
b[30618] == 30618 && 
b[30619] == 30619 && 
b[30620] == 30620 && 
b[30621] == 30621 && 
b[30622] == 30622 && 
b[30623] == 30623 && 
b[30624] == 30624 && 
b[30625] == 30625 && 
b[30626] == 30626 && 
b[30627] == 30627 && 
b[30628] == 30628 && 
b[30629] == 30629 && 
b[30630] == 30630 && 
b[30631] == 30631 && 
b[30632] == 30632 && 
b[30633] == 30633 && 
b[30634] == 30634 && 
b[30635] == 30635 && 
b[30636] == 30636 && 
b[30637] == 30637 && 
b[30638] == 30638 && 
b[30639] == 30639 && 
b[30640] == 30640 && 
b[30641] == 30641 && 
b[30642] == 30642 && 
b[30643] == 30643 && 
b[30644] == 30644 && 
b[30645] == 30645 && 
b[30646] == 30646 && 
b[30647] == 30647 && 
b[30648] == 30648 && 
b[30649] == 30649 && 
b[30650] == 30650 && 
b[30651] == 30651 && 
b[30652] == 30652 && 
b[30653] == 30653 && 
b[30654] == 30654 && 
b[30655] == 30655 && 
b[30656] == 30656 && 
b[30657] == 30657 && 
b[30658] == 30658 && 
b[30659] == 30659 && 
b[30660] == 30660 && 
b[30661] == 30661 && 
b[30662] == 30662 && 
b[30663] == 30663 && 
b[30664] == 30664 && 
b[30665] == 30665 && 
b[30666] == 30666 && 
b[30667] == 30667 && 
b[30668] == 30668 && 
b[30669] == 30669 && 
b[30670] == 30670 && 
b[30671] == 30671 && 
b[30672] == 30672 && 
b[30673] == 30673 && 
b[30674] == 30674 && 
b[30675] == 30675 && 
b[30676] == 30676 && 
b[30677] == 30677 && 
b[30678] == 30678 && 
b[30679] == 30679 && 
b[30680] == 30680 && 
b[30681] == 30681 && 
b[30682] == 30682 && 
b[30683] == 30683 && 
b[30684] == 30684 && 
b[30685] == 30685 && 
b[30686] == 30686 && 
b[30687] == 30687 && 
b[30688] == 30688 && 
b[30689] == 30689 && 
b[30690] == 30690 && 
b[30691] == 30691 && 
b[30692] == 30692 && 
b[30693] == 30693 && 
b[30694] == 30694 && 
b[30695] == 30695 && 
b[30696] == 30696 && 
b[30697] == 30697 && 
b[30698] == 30698 && 
b[30699] == 30699 && 
b[30700] == 30700 && 
b[30701] == 30701 && 
b[30702] == 30702 && 
b[30703] == 30703 && 
b[30704] == 30704 && 
b[30705] == 30705 && 
b[30706] == 30706 && 
b[30707] == 30707 && 
b[30708] == 30708 && 
b[30709] == 30709 && 
b[30710] == 30710 && 
b[30711] == 30711 && 
b[30712] == 30712 && 
b[30713] == 30713 && 
b[30714] == 30714 && 
b[30715] == 30715 && 
b[30716] == 30716 && 
b[30717] == 30717 && 
b[30718] == 30718 && 
b[30719] == 30719 && 
b[30720] == 30720 && 
b[30721] == 30721 && 
b[30722] == 30722 && 
b[30723] == 30723 && 
b[30724] == 30724 && 
b[30725] == 30725 && 
b[30726] == 30726 && 
b[30727] == 30727 && 
b[30728] == 30728 && 
b[30729] == 30729 && 
b[30730] == 30730 && 
b[30731] == 30731 && 
b[30732] == 30732 && 
b[30733] == 30733 && 
b[30734] == 30734 && 
b[30735] == 30735 && 
b[30736] == 30736 && 
b[30737] == 30737 && 
b[30738] == 30738 && 
b[30739] == 30739 && 
b[30740] == 30740 && 
b[30741] == 30741 && 
b[30742] == 30742 && 
b[30743] == 30743 && 
b[30744] == 30744 && 
b[30745] == 30745 && 
b[30746] == 30746 && 
b[30747] == 30747 && 
b[30748] == 30748 && 
b[30749] == 30749 && 
b[30750] == 30750 && 
b[30751] == 30751 && 
b[30752] == 30752 && 
b[30753] == 30753 && 
b[30754] == 30754 && 
b[30755] == 30755 && 
b[30756] == 30756 && 
b[30757] == 30757 && 
b[30758] == 30758 && 
b[30759] == 30759 && 
b[30760] == 30760 && 
b[30761] == 30761 && 
b[30762] == 30762 && 
b[30763] == 30763 && 
b[30764] == 30764 && 
b[30765] == 30765 && 
b[30766] == 30766 && 
b[30767] == 30767 && 
b[30768] == 30768 && 
b[30769] == 30769 && 
b[30770] == 30770 && 
b[30771] == 30771 && 
b[30772] == 30772 && 
b[30773] == 30773 && 
b[30774] == 30774 && 
b[30775] == 30775 && 
b[30776] == 30776 && 
b[30777] == 30777 && 
b[30778] == 30778 && 
b[30779] == 30779 && 
b[30780] == 30780 && 
b[30781] == 30781 && 
b[30782] == 30782 && 
b[30783] == 30783 && 
b[30784] == 30784 && 
b[30785] == 30785 && 
b[30786] == 30786 && 
b[30787] == 30787 && 
b[30788] == 30788 && 
b[30789] == 30789 && 
b[30790] == 30790 && 
b[30791] == 30791 && 
b[30792] == 30792 && 
b[30793] == 30793 && 
b[30794] == 30794 && 
b[30795] == 30795 && 
b[30796] == 30796 && 
b[30797] == 30797 && 
b[30798] == 30798 && 
b[30799] == 30799 && 
b[30800] == 30800 && 
b[30801] == 30801 && 
b[30802] == 30802 && 
b[30803] == 30803 && 
b[30804] == 30804 && 
b[30805] == 30805 && 
b[30806] == 30806 && 
b[30807] == 30807 && 
b[30808] == 30808 && 
b[30809] == 30809 && 
b[30810] == 30810 && 
b[30811] == 30811 && 
b[30812] == 30812 && 
b[30813] == 30813 && 
b[30814] == 30814 && 
b[30815] == 30815 && 
b[30816] == 30816 && 
b[30817] == 30817 && 
b[30818] == 30818 && 
b[30819] == 30819 && 
b[30820] == 30820 && 
b[30821] == 30821 && 
b[30822] == 30822 && 
b[30823] == 30823 && 
b[30824] == 30824 && 
b[30825] == 30825 && 
b[30826] == 30826 && 
b[30827] == 30827 && 
b[30828] == 30828 && 
b[30829] == 30829 && 
b[30830] == 30830 && 
b[30831] == 30831 && 
b[30832] == 30832 && 
b[30833] == 30833 && 
b[30834] == 30834 && 
b[30835] == 30835 && 
b[30836] == 30836 && 
b[30837] == 30837 && 
b[30838] == 30838 && 
b[30839] == 30839 && 
b[30840] == 30840 && 
b[30841] == 30841 && 
b[30842] == 30842 && 
b[30843] == 30843 && 
b[30844] == 30844 && 
b[30845] == 30845 && 
b[30846] == 30846 && 
b[30847] == 30847 && 
b[30848] == 30848 && 
b[30849] == 30849 && 
b[30850] == 30850 && 
b[30851] == 30851 && 
b[30852] == 30852 && 
b[30853] == 30853 && 
b[30854] == 30854 && 
b[30855] == 30855 && 
b[30856] == 30856 && 
b[30857] == 30857 && 
b[30858] == 30858 && 
b[30859] == 30859 && 
b[30860] == 30860 && 
b[30861] == 30861 && 
b[30862] == 30862 && 
b[30863] == 30863 && 
b[30864] == 30864 && 
b[30865] == 30865 && 
b[30866] == 30866 && 
b[30867] == 30867 && 
b[30868] == 30868 && 
b[30869] == 30869 && 
b[30870] == 30870 && 
b[30871] == 30871 && 
b[30872] == 30872 && 
b[30873] == 30873 && 
b[30874] == 30874 && 
b[30875] == 30875 && 
b[30876] == 30876 && 
b[30877] == 30877 && 
b[30878] == 30878 && 
b[30879] == 30879 && 
b[30880] == 30880 && 
b[30881] == 30881 && 
b[30882] == 30882 && 
b[30883] == 30883 && 
b[30884] == 30884 && 
b[30885] == 30885 && 
b[30886] == 30886 && 
b[30887] == 30887 && 
b[30888] == 30888 && 
b[30889] == 30889 && 
b[30890] == 30890 && 
b[30891] == 30891 && 
b[30892] == 30892 && 
b[30893] == 30893 && 
b[30894] == 30894 && 
b[30895] == 30895 && 
b[30896] == 30896 && 
b[30897] == 30897 && 
b[30898] == 30898 && 
b[30899] == 30899 && 
b[30900] == 30900 && 
b[30901] == 30901 && 
b[30902] == 30902 && 
b[30903] == 30903 && 
b[30904] == 30904 && 
b[30905] == 30905 && 
b[30906] == 30906 && 
b[30907] == 30907 && 
b[30908] == 30908 && 
b[30909] == 30909 && 
b[30910] == 30910 && 
b[30911] == 30911 && 
b[30912] == 30912 && 
b[30913] == 30913 && 
b[30914] == 30914 && 
b[30915] == 30915 && 
b[30916] == 30916 && 
b[30917] == 30917 && 
b[30918] == 30918 && 
b[30919] == 30919 && 
b[30920] == 30920 && 
b[30921] == 30921 && 
b[30922] == 30922 && 
b[30923] == 30923 && 
b[30924] == 30924 && 
b[30925] == 30925 && 
b[30926] == 30926 && 
b[30927] == 30927 && 
b[30928] == 30928 && 
b[30929] == 30929 && 
b[30930] == 30930 && 
b[30931] == 30931 && 
b[30932] == 30932 && 
b[30933] == 30933 && 
b[30934] == 30934 && 
b[30935] == 30935 && 
b[30936] == 30936 && 
b[30937] == 30937 && 
b[30938] == 30938 && 
b[30939] == 30939 && 
b[30940] == 30940 && 
b[30941] == 30941 && 
b[30942] == 30942 && 
b[30943] == 30943 && 
b[30944] == 30944 && 
b[30945] == 30945 && 
b[30946] == 30946 && 
b[30947] == 30947 && 
b[30948] == 30948 && 
b[30949] == 30949 && 
b[30950] == 30950 && 
b[30951] == 30951 && 
b[30952] == 30952 && 
b[30953] == 30953 && 
b[30954] == 30954 && 
b[30955] == 30955 && 
b[30956] == 30956 && 
b[30957] == 30957 && 
b[30958] == 30958 && 
b[30959] == 30959 && 
b[30960] == 30960 && 
b[30961] == 30961 && 
b[30962] == 30962 && 
b[30963] == 30963 && 
b[30964] == 30964 && 
b[30965] == 30965 && 
b[30966] == 30966 && 
b[30967] == 30967 && 
b[30968] == 30968 && 
b[30969] == 30969 && 
b[30970] == 30970 && 
b[30971] == 30971 && 
b[30972] == 30972 && 
b[30973] == 30973 && 
b[30974] == 30974 && 
b[30975] == 30975 && 
b[30976] == 30976 && 
b[30977] == 30977 && 
b[30978] == 30978 && 
b[30979] == 30979 && 
b[30980] == 30980 && 
b[30981] == 30981 && 
b[30982] == 30982 && 
b[30983] == 30983 && 
b[30984] == 30984 && 
b[30985] == 30985 && 
b[30986] == 30986 && 
b[30987] == 30987 && 
b[30988] == 30988 && 
b[30989] == 30989 && 
b[30990] == 30990 && 
b[30991] == 30991 && 
b[30992] == 30992 && 
b[30993] == 30993 && 
b[30994] == 30994 && 
b[30995] == 30995 && 
b[30996] == 30996 && 
b[30997] == 30997 && 
b[30998] == 30998 && 
b[30999] == 30999 && 
b[31000] == 31000 && 
b[31001] == 31001 && 
b[31002] == 31002 && 
b[31003] == 31003 && 
b[31004] == 31004 && 
b[31005] == 31005 && 
b[31006] == 31006 && 
b[31007] == 31007 && 
b[31008] == 31008 && 
b[31009] == 31009 && 
b[31010] == 31010 && 
b[31011] == 31011 && 
b[31012] == 31012 && 
b[31013] == 31013 && 
b[31014] == 31014 && 
b[31015] == 31015 && 
b[31016] == 31016 && 
b[31017] == 31017 && 
b[31018] == 31018 && 
b[31019] == 31019 && 
b[31020] == 31020 && 
b[31021] == 31021 && 
b[31022] == 31022 && 
b[31023] == 31023 && 
b[31024] == 31024 && 
b[31025] == 31025 && 
b[31026] == 31026 && 
b[31027] == 31027 && 
b[31028] == 31028 && 
b[31029] == 31029 && 
b[31030] == 31030 && 
b[31031] == 31031 && 
b[31032] == 31032 && 
b[31033] == 31033 && 
b[31034] == 31034 && 
b[31035] == 31035 && 
b[31036] == 31036 && 
b[31037] == 31037 && 
b[31038] == 31038 && 
b[31039] == 31039 && 
b[31040] == 31040 && 
b[31041] == 31041 && 
b[31042] == 31042 && 
b[31043] == 31043 && 
b[31044] == 31044 && 
b[31045] == 31045 && 
b[31046] == 31046 && 
b[31047] == 31047 && 
b[31048] == 31048 && 
b[31049] == 31049 && 
b[31050] == 31050 && 
b[31051] == 31051 && 
b[31052] == 31052 && 
b[31053] == 31053 && 
b[31054] == 31054 && 
b[31055] == 31055 && 
b[31056] == 31056 && 
b[31057] == 31057 && 
b[31058] == 31058 && 
b[31059] == 31059 && 
b[31060] == 31060 && 
b[31061] == 31061 && 
b[31062] == 31062 && 
b[31063] == 31063 && 
b[31064] == 31064 && 
b[31065] == 31065 && 
b[31066] == 31066 && 
b[31067] == 31067 && 
b[31068] == 31068 && 
b[31069] == 31069 && 
b[31070] == 31070 && 
b[31071] == 31071 && 
b[31072] == 31072 && 
b[31073] == 31073 && 
b[31074] == 31074 && 
b[31075] == 31075 && 
b[31076] == 31076 && 
b[31077] == 31077 && 
b[31078] == 31078 && 
b[31079] == 31079 && 
b[31080] == 31080 && 
b[31081] == 31081 && 
b[31082] == 31082 && 
b[31083] == 31083 && 
b[31084] == 31084 && 
b[31085] == 31085 && 
b[31086] == 31086 && 
b[31087] == 31087 && 
b[31088] == 31088 && 
b[31089] == 31089 && 
b[31090] == 31090 && 
b[31091] == 31091 && 
b[31092] == 31092 && 
b[31093] == 31093 && 
b[31094] == 31094 && 
b[31095] == 31095 && 
b[31096] == 31096 && 
b[31097] == 31097 && 
b[31098] == 31098 && 
b[31099] == 31099 && 
b[31100] == 31100 && 
b[31101] == 31101 && 
b[31102] == 31102 && 
b[31103] == 31103 && 
b[31104] == 31104 && 
b[31105] == 31105 && 
b[31106] == 31106 && 
b[31107] == 31107 && 
b[31108] == 31108 && 
b[31109] == 31109 && 
b[31110] == 31110 && 
b[31111] == 31111 && 
b[31112] == 31112 && 
b[31113] == 31113 && 
b[31114] == 31114 && 
b[31115] == 31115 && 
b[31116] == 31116 && 
b[31117] == 31117 && 
b[31118] == 31118 && 
b[31119] == 31119 && 
b[31120] == 31120 && 
b[31121] == 31121 && 
b[31122] == 31122 && 
b[31123] == 31123 && 
b[31124] == 31124 && 
b[31125] == 31125 && 
b[31126] == 31126 && 
b[31127] == 31127 && 
b[31128] == 31128 && 
b[31129] == 31129 && 
b[31130] == 31130 && 
b[31131] == 31131 && 
b[31132] == 31132 && 
b[31133] == 31133 && 
b[31134] == 31134 && 
b[31135] == 31135 && 
b[31136] == 31136 && 
b[31137] == 31137 && 
b[31138] == 31138 && 
b[31139] == 31139 && 
b[31140] == 31140 && 
b[31141] == 31141 && 
b[31142] == 31142 && 
b[31143] == 31143 && 
b[31144] == 31144 && 
b[31145] == 31145 && 
b[31146] == 31146 && 
b[31147] == 31147 && 
b[31148] == 31148 && 
b[31149] == 31149 && 
b[31150] == 31150 && 
b[31151] == 31151 && 
b[31152] == 31152 && 
b[31153] == 31153 && 
b[31154] == 31154 && 
b[31155] == 31155 && 
b[31156] == 31156 && 
b[31157] == 31157 && 
b[31158] == 31158 && 
b[31159] == 31159 && 
b[31160] == 31160 && 
b[31161] == 31161 && 
b[31162] == 31162 && 
b[31163] == 31163 && 
b[31164] == 31164 && 
b[31165] == 31165 && 
b[31166] == 31166 && 
b[31167] == 31167 && 
b[31168] == 31168 && 
b[31169] == 31169 && 
b[31170] == 31170 && 
b[31171] == 31171 && 
b[31172] == 31172 && 
b[31173] == 31173 && 
b[31174] == 31174 && 
b[31175] == 31175 && 
b[31176] == 31176 && 
b[31177] == 31177 && 
b[31178] == 31178 && 
b[31179] == 31179 && 
b[31180] == 31180 && 
b[31181] == 31181 && 
b[31182] == 31182 && 
b[31183] == 31183 && 
b[31184] == 31184 && 
b[31185] == 31185 && 
b[31186] == 31186 && 
b[31187] == 31187 && 
b[31188] == 31188 && 
b[31189] == 31189 && 
b[31190] == 31190 && 
b[31191] == 31191 && 
b[31192] == 31192 && 
b[31193] == 31193 && 
b[31194] == 31194 && 
b[31195] == 31195 && 
b[31196] == 31196 && 
b[31197] == 31197 && 
b[31198] == 31198 && 
b[31199] == 31199 && 
b[31200] == 31200 && 
b[31201] == 31201 && 
b[31202] == 31202 && 
b[31203] == 31203 && 
b[31204] == 31204 && 
b[31205] == 31205 && 
b[31206] == 31206 && 
b[31207] == 31207 && 
b[31208] == 31208 && 
b[31209] == 31209 && 
b[31210] == 31210 && 
b[31211] == 31211 && 
b[31212] == 31212 && 
b[31213] == 31213 && 
b[31214] == 31214 && 
b[31215] == 31215 && 
b[31216] == 31216 && 
b[31217] == 31217 && 
b[31218] == 31218 && 
b[31219] == 31219 && 
b[31220] == 31220 && 
b[31221] == 31221 && 
b[31222] == 31222 && 
b[31223] == 31223 && 
b[31224] == 31224 && 
b[31225] == 31225 && 
b[31226] == 31226 && 
b[31227] == 31227 && 
b[31228] == 31228 && 
b[31229] == 31229 && 
b[31230] == 31230 && 
b[31231] == 31231 && 
b[31232] == 31232 && 
b[31233] == 31233 && 
b[31234] == 31234 && 
b[31235] == 31235 && 
b[31236] == 31236 && 
b[31237] == 31237 && 
b[31238] == 31238 && 
b[31239] == 31239 && 
b[31240] == 31240 && 
b[31241] == 31241 && 
b[31242] == 31242 && 
b[31243] == 31243 && 
b[31244] == 31244 && 
b[31245] == 31245 && 
b[31246] == 31246 && 
b[31247] == 31247 && 
b[31248] == 31248 && 
b[31249] == 31249 && 
b[31250] == 31250 && 
b[31251] == 31251 && 
b[31252] == 31252 && 
b[31253] == 31253 && 
b[31254] == 31254 && 
b[31255] == 31255 && 
b[31256] == 31256 && 
b[31257] == 31257 && 
b[31258] == 31258 && 
b[31259] == 31259 && 
b[31260] == 31260 && 
b[31261] == 31261 && 
b[31262] == 31262 && 
b[31263] == 31263 && 
b[31264] == 31264 && 
b[31265] == 31265 && 
b[31266] == 31266 && 
b[31267] == 31267 && 
b[31268] == 31268 && 
b[31269] == 31269 && 
b[31270] == 31270 && 
b[31271] == 31271 && 
b[31272] == 31272 && 
b[31273] == 31273 && 
b[31274] == 31274 && 
b[31275] == 31275 && 
b[31276] == 31276 && 
b[31277] == 31277 && 
b[31278] == 31278 && 
b[31279] == 31279 && 
b[31280] == 31280 && 
b[31281] == 31281 && 
b[31282] == 31282 && 
b[31283] == 31283 && 
b[31284] == 31284 && 
b[31285] == 31285 && 
b[31286] == 31286 && 
b[31287] == 31287 && 
b[31288] == 31288 && 
b[31289] == 31289 && 
b[31290] == 31290 && 
b[31291] == 31291 && 
b[31292] == 31292 && 
b[31293] == 31293 && 
b[31294] == 31294 && 
b[31295] == 31295 && 
b[31296] == 31296 && 
b[31297] == 31297 && 
b[31298] == 31298 && 
b[31299] == 31299 && 
b[31300] == 31300 && 
b[31301] == 31301 && 
b[31302] == 31302 && 
b[31303] == 31303 && 
b[31304] == 31304 && 
b[31305] == 31305 && 
b[31306] == 31306 && 
b[31307] == 31307 && 
b[31308] == 31308 && 
b[31309] == 31309 && 
b[31310] == 31310 && 
b[31311] == 31311 && 
b[31312] == 31312 && 
b[31313] == 31313 && 
b[31314] == 31314 && 
b[31315] == 31315 && 
b[31316] == 31316 && 
b[31317] == 31317 && 
b[31318] == 31318 && 
b[31319] == 31319 && 
b[31320] == 31320 && 
b[31321] == 31321 && 
b[31322] == 31322 && 
b[31323] == 31323 && 
b[31324] == 31324 && 
b[31325] == 31325 && 
b[31326] == 31326 && 
b[31327] == 31327 && 
b[31328] == 31328 && 
b[31329] == 31329 && 
b[31330] == 31330 && 
b[31331] == 31331 && 
b[31332] == 31332 && 
b[31333] == 31333 && 
b[31334] == 31334 && 
b[31335] == 31335 && 
b[31336] == 31336 && 
b[31337] == 31337 && 
b[31338] == 31338 && 
b[31339] == 31339 && 
b[31340] == 31340 && 
b[31341] == 31341 && 
b[31342] == 31342 && 
b[31343] == 31343 && 
b[31344] == 31344 && 
b[31345] == 31345 && 
b[31346] == 31346 && 
b[31347] == 31347 && 
b[31348] == 31348 && 
b[31349] == 31349 && 
b[31350] == 31350 && 
b[31351] == 31351 && 
b[31352] == 31352 && 
b[31353] == 31353 && 
b[31354] == 31354 && 
b[31355] == 31355 && 
b[31356] == 31356 && 
b[31357] == 31357 && 
b[31358] == 31358 && 
b[31359] == 31359 && 
b[31360] == 31360 && 
b[31361] == 31361 && 
b[31362] == 31362 && 
b[31363] == 31363 && 
b[31364] == 31364 && 
b[31365] == 31365 && 
b[31366] == 31366 && 
b[31367] == 31367 && 
b[31368] == 31368 && 
b[31369] == 31369 && 
b[31370] == 31370 && 
b[31371] == 31371 && 
b[31372] == 31372 && 
b[31373] == 31373 && 
b[31374] == 31374 && 
b[31375] == 31375 && 
b[31376] == 31376 && 
b[31377] == 31377 && 
b[31378] == 31378 && 
b[31379] == 31379 && 
b[31380] == 31380 && 
b[31381] == 31381 && 
b[31382] == 31382 && 
b[31383] == 31383 && 
b[31384] == 31384 && 
b[31385] == 31385 && 
b[31386] == 31386 && 
b[31387] == 31387 && 
b[31388] == 31388 && 
b[31389] == 31389 && 
b[31390] == 31390 && 
b[31391] == 31391 && 
b[31392] == 31392 && 
b[31393] == 31393 && 
b[31394] == 31394 && 
b[31395] == 31395 && 
b[31396] == 31396 && 
b[31397] == 31397 && 
b[31398] == 31398 && 
b[31399] == 31399 && 
b[31400] == 31400 && 
b[31401] == 31401 && 
b[31402] == 31402 && 
b[31403] == 31403 && 
b[31404] == 31404 && 
b[31405] == 31405 && 
b[31406] == 31406 && 
b[31407] == 31407 && 
b[31408] == 31408 && 
b[31409] == 31409 && 
b[31410] == 31410 && 
b[31411] == 31411 && 
b[31412] == 31412 && 
b[31413] == 31413 && 
b[31414] == 31414 && 
b[31415] == 31415 && 
b[31416] == 31416 && 
b[31417] == 31417 && 
b[31418] == 31418 && 
b[31419] == 31419 && 
b[31420] == 31420 && 
b[31421] == 31421 && 
b[31422] == 31422 && 
b[31423] == 31423 && 
b[31424] == 31424 && 
b[31425] == 31425 && 
b[31426] == 31426 && 
b[31427] == 31427 && 
b[31428] == 31428 && 
b[31429] == 31429 && 
b[31430] == 31430 && 
b[31431] == 31431 && 
b[31432] == 31432 && 
b[31433] == 31433 && 
b[31434] == 31434 && 
b[31435] == 31435 && 
b[31436] == 31436 && 
b[31437] == 31437 && 
b[31438] == 31438 && 
b[31439] == 31439 && 
b[31440] == 31440 && 
b[31441] == 31441 && 
b[31442] == 31442 && 
b[31443] == 31443 && 
b[31444] == 31444 && 
b[31445] == 31445 && 
b[31446] == 31446 && 
b[31447] == 31447 && 
b[31448] == 31448 && 
b[31449] == 31449 && 
b[31450] == 31450 && 
b[31451] == 31451 && 
b[31452] == 31452 && 
b[31453] == 31453 && 
b[31454] == 31454 && 
b[31455] == 31455 && 
b[31456] == 31456 && 
b[31457] == 31457 && 
b[31458] == 31458 && 
b[31459] == 31459 && 
b[31460] == 31460 && 
b[31461] == 31461 && 
b[31462] == 31462 && 
b[31463] == 31463 && 
b[31464] == 31464 && 
b[31465] == 31465 && 
b[31466] == 31466 && 
b[31467] == 31467 && 
b[31468] == 31468 && 
b[31469] == 31469 && 
b[31470] == 31470 && 
b[31471] == 31471 && 
b[31472] == 31472 && 
b[31473] == 31473 && 
b[31474] == 31474 && 
b[31475] == 31475 && 
b[31476] == 31476 && 
b[31477] == 31477 && 
b[31478] == 31478 && 
b[31479] == 31479 && 
b[31480] == 31480 && 
b[31481] == 31481 && 
b[31482] == 31482 && 
b[31483] == 31483 && 
b[31484] == 31484 && 
b[31485] == 31485 && 
b[31486] == 31486 && 
b[31487] == 31487 && 
b[31488] == 31488 && 
b[31489] == 31489 && 
b[31490] == 31490 && 
b[31491] == 31491 && 
b[31492] == 31492 && 
b[31493] == 31493 && 
b[31494] == 31494 && 
b[31495] == 31495 && 
b[31496] == 31496 && 
b[31497] == 31497 && 
b[31498] == 31498 && 
b[31499] == 31499 && 
b[31500] == 31500 && 
b[31501] == 31501 && 
b[31502] == 31502 && 
b[31503] == 31503 && 
b[31504] == 31504 && 
b[31505] == 31505 && 
b[31506] == 31506 && 
b[31507] == 31507 && 
b[31508] == 31508 && 
b[31509] == 31509 && 
b[31510] == 31510 && 
b[31511] == 31511 && 
b[31512] == 31512 && 
b[31513] == 31513 && 
b[31514] == 31514 && 
b[31515] == 31515 && 
b[31516] == 31516 && 
b[31517] == 31517 && 
b[31518] == 31518 && 
b[31519] == 31519 && 
b[31520] == 31520 && 
b[31521] == 31521 && 
b[31522] == 31522 && 
b[31523] == 31523 && 
b[31524] == 31524 && 
b[31525] == 31525 && 
b[31526] == 31526 && 
b[31527] == 31527 && 
b[31528] == 31528 && 
b[31529] == 31529 && 
b[31530] == 31530 && 
b[31531] == 31531 && 
b[31532] == 31532 && 
b[31533] == 31533 && 
b[31534] == 31534 && 
b[31535] == 31535 && 
b[31536] == 31536 && 
b[31537] == 31537 && 
b[31538] == 31538 && 
b[31539] == 31539 && 
b[31540] == 31540 && 
b[31541] == 31541 && 
b[31542] == 31542 && 
b[31543] == 31543 && 
b[31544] == 31544 && 
b[31545] == 31545 && 
b[31546] == 31546 && 
b[31547] == 31547 && 
b[31548] == 31548 && 
b[31549] == 31549 && 
b[31550] == 31550 && 
b[31551] == 31551 && 
b[31552] == 31552 && 
b[31553] == 31553 && 
b[31554] == 31554 && 
b[31555] == 31555 && 
b[31556] == 31556 && 
b[31557] == 31557 && 
b[31558] == 31558 && 
b[31559] == 31559 && 
b[31560] == 31560 && 
b[31561] == 31561 && 
b[31562] == 31562 && 
b[31563] == 31563 && 
b[31564] == 31564 && 
b[31565] == 31565 && 
b[31566] == 31566 && 
b[31567] == 31567 && 
b[31568] == 31568 && 
b[31569] == 31569 && 
b[31570] == 31570 && 
b[31571] == 31571 && 
b[31572] == 31572 && 
b[31573] == 31573 && 
b[31574] == 31574 && 
b[31575] == 31575 && 
b[31576] == 31576 && 
b[31577] == 31577 && 
b[31578] == 31578 && 
b[31579] == 31579 && 
b[31580] == 31580 && 
b[31581] == 31581 && 
b[31582] == 31582 && 
b[31583] == 31583 && 
b[31584] == 31584 && 
b[31585] == 31585 && 
b[31586] == 31586 && 
b[31587] == 31587 && 
b[31588] == 31588 && 
b[31589] == 31589 && 
b[31590] == 31590 && 
b[31591] == 31591 && 
b[31592] == 31592 && 
b[31593] == 31593 && 
b[31594] == 31594 && 
b[31595] == 31595 && 
b[31596] == 31596 && 
b[31597] == 31597 && 
b[31598] == 31598 && 
b[31599] == 31599 && 
b[31600] == 31600 && 
b[31601] == 31601 && 
b[31602] == 31602 && 
b[31603] == 31603 && 
b[31604] == 31604 && 
b[31605] == 31605 && 
b[31606] == 31606 && 
b[31607] == 31607 && 
b[31608] == 31608 && 
b[31609] == 31609 && 
b[31610] == 31610 && 
b[31611] == 31611 && 
b[31612] == 31612 && 
b[31613] == 31613 && 
b[31614] == 31614 && 
b[31615] == 31615 && 
b[31616] == 31616 && 
b[31617] == 31617 && 
b[31618] == 31618 && 
b[31619] == 31619 && 
b[31620] == 31620 && 
b[31621] == 31621 && 
b[31622] == 31622 && 
b[31623] == 31623 && 
b[31624] == 31624 && 
b[31625] == 31625 && 
b[31626] == 31626 && 
b[31627] == 31627 && 
b[31628] == 31628 && 
b[31629] == 31629 && 
b[31630] == 31630 && 
b[31631] == 31631 && 
b[31632] == 31632 && 
b[31633] == 31633 && 
b[31634] == 31634 && 
b[31635] == 31635 && 
b[31636] == 31636 && 
b[31637] == 31637 && 
b[31638] == 31638 && 
b[31639] == 31639 && 
b[31640] == 31640 && 
b[31641] == 31641 && 
b[31642] == 31642 && 
b[31643] == 31643 && 
b[31644] == 31644 && 
b[31645] == 31645 && 
b[31646] == 31646 && 
b[31647] == 31647 && 
b[31648] == 31648 && 
b[31649] == 31649 && 
b[31650] == 31650 && 
b[31651] == 31651 && 
b[31652] == 31652 && 
b[31653] == 31653 && 
b[31654] == 31654 && 
b[31655] == 31655 && 
b[31656] == 31656 && 
b[31657] == 31657 && 
b[31658] == 31658 && 
b[31659] == 31659 && 
b[31660] == 31660 && 
b[31661] == 31661 && 
b[31662] == 31662 && 
b[31663] == 31663 && 
b[31664] == 31664 && 
b[31665] == 31665 && 
b[31666] == 31666 && 
b[31667] == 31667 && 
b[31668] == 31668 && 
b[31669] == 31669 && 
b[31670] == 31670 && 
b[31671] == 31671 && 
b[31672] == 31672 && 
b[31673] == 31673 && 
b[31674] == 31674 && 
b[31675] == 31675 && 
b[31676] == 31676 && 
b[31677] == 31677 && 
b[31678] == 31678 && 
b[31679] == 31679 && 
b[31680] == 31680 && 
b[31681] == 31681 && 
b[31682] == 31682 && 
b[31683] == 31683 && 
b[31684] == 31684 && 
b[31685] == 31685 && 
b[31686] == 31686 && 
b[31687] == 31687 && 
b[31688] == 31688 && 
b[31689] == 31689 && 
b[31690] == 31690 && 
b[31691] == 31691 && 
b[31692] == 31692 && 
b[31693] == 31693 && 
b[31694] == 31694 && 
b[31695] == 31695 && 
b[31696] == 31696 && 
b[31697] == 31697 && 
b[31698] == 31698 && 
b[31699] == 31699 && 
b[31700] == 31700 && 
b[31701] == 31701 && 
b[31702] == 31702 && 
b[31703] == 31703 && 
b[31704] == 31704 && 
b[31705] == 31705 && 
b[31706] == 31706 && 
b[31707] == 31707 && 
b[31708] == 31708 && 
b[31709] == 31709 && 
b[31710] == 31710 && 
b[31711] == 31711 && 
b[31712] == 31712 && 
b[31713] == 31713 && 
b[31714] == 31714 && 
b[31715] == 31715 && 
b[31716] == 31716 && 
b[31717] == 31717 && 
b[31718] == 31718 && 
b[31719] == 31719 && 
b[31720] == 31720 && 
b[31721] == 31721 && 
b[31722] == 31722 && 
b[31723] == 31723 && 
b[31724] == 31724 && 
b[31725] == 31725 && 
b[31726] == 31726 && 
b[31727] == 31727 && 
b[31728] == 31728 && 
b[31729] == 31729 && 
b[31730] == 31730 && 
b[31731] == 31731 && 
b[31732] == 31732 && 
b[31733] == 31733 && 
b[31734] == 31734 && 
b[31735] == 31735 && 
b[31736] == 31736 && 
b[31737] == 31737 && 
b[31738] == 31738 && 
b[31739] == 31739 && 
b[31740] == 31740 && 
b[31741] == 31741 && 
b[31742] == 31742 && 
b[31743] == 31743 && 
b[31744] == 31744 && 
b[31745] == 31745 && 
b[31746] == 31746 && 
b[31747] == 31747 && 
b[31748] == 31748 && 
b[31749] == 31749 && 
b[31750] == 31750 && 
b[31751] == 31751 && 
b[31752] == 31752 && 
b[31753] == 31753 && 
b[31754] == 31754 && 
b[31755] == 31755 && 
b[31756] == 31756 && 
b[31757] == 31757 && 
b[31758] == 31758 && 
b[31759] == 31759 && 
b[31760] == 31760 && 
b[31761] == 31761 && 
b[31762] == 31762 && 
b[31763] == 31763 && 
b[31764] == 31764 && 
b[31765] == 31765 && 
b[31766] == 31766 && 
b[31767] == 31767 && 
b[31768] == 31768 && 
b[31769] == 31769 && 
b[31770] == 31770 && 
b[31771] == 31771 && 
b[31772] == 31772 && 
b[31773] == 31773 && 
b[31774] == 31774 && 
b[31775] == 31775 && 
b[31776] == 31776 && 
b[31777] == 31777 && 
b[31778] == 31778 && 
b[31779] == 31779 && 
b[31780] == 31780 && 
b[31781] == 31781 && 
b[31782] == 31782 && 
b[31783] == 31783 && 
b[31784] == 31784 && 
b[31785] == 31785 && 
b[31786] == 31786 && 
b[31787] == 31787 && 
b[31788] == 31788 && 
b[31789] == 31789 && 
b[31790] == 31790 && 
b[31791] == 31791 && 
b[31792] == 31792 && 
b[31793] == 31793 && 
b[31794] == 31794 && 
b[31795] == 31795 && 
b[31796] == 31796 && 
b[31797] == 31797 && 
b[31798] == 31798 && 
b[31799] == 31799 && 
b[31800] == 31800 && 
b[31801] == 31801 && 
b[31802] == 31802 && 
b[31803] == 31803 && 
b[31804] == 31804 && 
b[31805] == 31805 && 
b[31806] == 31806 && 
b[31807] == 31807 && 
b[31808] == 31808 && 
b[31809] == 31809 && 
b[31810] == 31810 && 
b[31811] == 31811 && 
b[31812] == 31812 && 
b[31813] == 31813 && 
b[31814] == 31814 && 
b[31815] == 31815 && 
b[31816] == 31816 && 
b[31817] == 31817 && 
b[31818] == 31818 && 
b[31819] == 31819 && 
b[31820] == 31820 && 
b[31821] == 31821 && 
b[31822] == 31822 && 
b[31823] == 31823 && 
b[31824] == 31824 && 
b[31825] == 31825 && 
b[31826] == 31826 && 
b[31827] == 31827 && 
b[31828] == 31828 && 
b[31829] == 31829 && 
b[31830] == 31830 && 
b[31831] == 31831 && 
b[31832] == 31832 && 
b[31833] == 31833 && 
b[31834] == 31834 && 
b[31835] == 31835 && 
b[31836] == 31836 && 
b[31837] == 31837 && 
b[31838] == 31838 && 
b[31839] == 31839 && 
b[31840] == 31840 && 
b[31841] == 31841 && 
b[31842] == 31842 && 
b[31843] == 31843 && 
b[31844] == 31844 && 
b[31845] == 31845 && 
b[31846] == 31846 && 
b[31847] == 31847 && 
b[31848] == 31848 && 
b[31849] == 31849 && 
b[31850] == 31850 && 
b[31851] == 31851 && 
b[31852] == 31852 && 
b[31853] == 31853 && 
b[31854] == 31854 && 
b[31855] == 31855 && 
b[31856] == 31856 && 
b[31857] == 31857 && 
b[31858] == 31858 && 
b[31859] == 31859 && 
b[31860] == 31860 && 
b[31861] == 31861 && 
b[31862] == 31862 && 
b[31863] == 31863 && 
b[31864] == 31864 && 
b[31865] == 31865 && 
b[31866] == 31866 && 
b[31867] == 31867 && 
b[31868] == 31868 && 
b[31869] == 31869 && 
b[31870] == 31870 && 
b[31871] == 31871 && 
b[31872] == 31872 && 
b[31873] == 31873 && 
b[31874] == 31874 && 
b[31875] == 31875 && 
b[31876] == 31876 && 
b[31877] == 31877 && 
b[31878] == 31878 && 
b[31879] == 31879 && 
b[31880] == 31880 && 
b[31881] == 31881 && 
b[31882] == 31882 && 
b[31883] == 31883 && 
b[31884] == 31884 && 
b[31885] == 31885 && 
b[31886] == 31886 && 
b[31887] == 31887 && 
b[31888] == 31888 && 
b[31889] == 31889 && 
b[31890] == 31890 && 
b[31891] == 31891 && 
b[31892] == 31892 && 
b[31893] == 31893 && 
b[31894] == 31894 && 
b[31895] == 31895 && 
b[31896] == 31896 && 
b[31897] == 31897 && 
b[31898] == 31898 && 
b[31899] == 31899 && 
b[31900] == 31900 && 
b[31901] == 31901 && 
b[31902] == 31902 && 
b[31903] == 31903 && 
b[31904] == 31904 && 
b[31905] == 31905 && 
b[31906] == 31906 && 
b[31907] == 31907 && 
b[31908] == 31908 && 
b[31909] == 31909 && 
b[31910] == 31910 && 
b[31911] == 31911 && 
b[31912] == 31912 && 
b[31913] == 31913 && 
b[31914] == 31914 && 
b[31915] == 31915 && 
b[31916] == 31916 && 
b[31917] == 31917 && 
b[31918] == 31918 && 
b[31919] == 31919 && 
b[31920] == 31920 && 
b[31921] == 31921 && 
b[31922] == 31922 && 
b[31923] == 31923 && 
b[31924] == 31924 && 
b[31925] == 31925 && 
b[31926] == 31926 && 
b[31927] == 31927 && 
b[31928] == 31928 && 
b[31929] == 31929 && 
b[31930] == 31930 && 
b[31931] == 31931 && 
b[31932] == 31932 && 
b[31933] == 31933 && 
b[31934] == 31934 && 
b[31935] == 31935 && 
b[31936] == 31936 && 
b[31937] == 31937 && 
b[31938] == 31938 && 
b[31939] == 31939 && 
b[31940] == 31940 && 
b[31941] == 31941 && 
b[31942] == 31942 && 
b[31943] == 31943 && 
b[31944] == 31944 && 
b[31945] == 31945 && 
b[31946] == 31946 && 
b[31947] == 31947 && 
b[31948] == 31948 && 
b[31949] == 31949 && 
b[31950] == 31950 && 
b[31951] == 31951 && 
b[31952] == 31952 && 
b[31953] == 31953 && 
b[31954] == 31954 && 
b[31955] == 31955 && 
b[31956] == 31956 && 
b[31957] == 31957 && 
b[31958] == 31958 && 
b[31959] == 31959 && 
b[31960] == 31960 && 
b[31961] == 31961 && 
b[31962] == 31962 && 
b[31963] == 31963 && 
b[31964] == 31964 && 
b[31965] == 31965 && 
b[31966] == 31966 && 
b[31967] == 31967 && 
b[31968] == 31968 && 
b[31969] == 31969 && 
b[31970] == 31970 && 
b[31971] == 31971 && 
b[31972] == 31972 && 
b[31973] == 31973 && 
b[31974] == 31974 && 
b[31975] == 31975 && 
b[31976] == 31976 && 
b[31977] == 31977 && 
b[31978] == 31978 && 
b[31979] == 31979 && 
b[31980] == 31980 && 
b[31981] == 31981 && 
b[31982] == 31982 && 
b[31983] == 31983 && 
b[31984] == 31984 && 
b[31985] == 31985 && 
b[31986] == 31986 && 
b[31987] == 31987 && 
b[31988] == 31988 && 
b[31989] == 31989 && 
b[31990] == 31990 && 
b[31991] == 31991 && 
b[31992] == 31992 && 
b[31993] == 31993 && 
b[31994] == 31994 && 
b[31995] == 31995 && 
b[31996] == 31996 && 
b[31997] == 31997 && 
b[31998] == 31998 && 
b[31999] == 31999 && 
b[32000] == 32000 && 
b[32001] == 32001 && 
b[32002] == 32002 && 
b[32003] == 32003 && 
b[32004] == 32004 && 
b[32005] == 32005 && 
b[32006] == 32006 && 
b[32007] == 32007 && 
b[32008] == 32008 && 
b[32009] == 32009 && 
b[32010] == 32010 && 
b[32011] == 32011 && 
b[32012] == 32012 && 
b[32013] == 32013 && 
b[32014] == 32014 && 
b[32015] == 32015 && 
b[32016] == 32016 && 
b[32017] == 32017 && 
b[32018] == 32018 && 
b[32019] == 32019 && 
b[32020] == 32020 && 
b[32021] == 32021 && 
b[32022] == 32022 && 
b[32023] == 32023 && 
b[32024] == 32024 && 
b[32025] == 32025 && 
b[32026] == 32026 && 
b[32027] == 32027 && 
b[32028] == 32028 && 
b[32029] == 32029 && 
b[32030] == 32030 && 
b[32031] == 32031 && 
b[32032] == 32032 && 
b[32033] == 32033 && 
b[32034] == 32034 && 
b[32035] == 32035 && 
b[32036] == 32036 && 
b[32037] == 32037 && 
b[32038] == 32038 && 
b[32039] == 32039 && 
b[32040] == 32040 && 
b[32041] == 32041 && 
b[32042] == 32042 && 
b[32043] == 32043 && 
b[32044] == 32044 && 
b[32045] == 32045 && 
b[32046] == 32046 && 
b[32047] == 32047 && 
b[32048] == 32048 && 
b[32049] == 32049 && 
b[32050] == 32050 && 
b[32051] == 32051 && 
b[32052] == 32052 && 
b[32053] == 32053 && 
b[32054] == 32054 && 
b[32055] == 32055 && 
b[32056] == 32056 && 
b[32057] == 32057 && 
b[32058] == 32058 && 
b[32059] == 32059 && 
b[32060] == 32060 && 
b[32061] == 32061 && 
b[32062] == 32062 && 
b[32063] == 32063 && 
b[32064] == 32064 && 
b[32065] == 32065 && 
b[32066] == 32066 && 
b[32067] == 32067 && 
b[32068] == 32068 && 
b[32069] == 32069 && 
b[32070] == 32070 && 
b[32071] == 32071 && 
b[32072] == 32072 && 
b[32073] == 32073 && 
b[32074] == 32074 && 
b[32075] == 32075 && 
b[32076] == 32076 && 
b[32077] == 32077 && 
b[32078] == 32078 && 
b[32079] == 32079 && 
b[32080] == 32080 && 
b[32081] == 32081 && 
b[32082] == 32082 && 
b[32083] == 32083 && 
b[32084] == 32084 && 
b[32085] == 32085 && 
b[32086] == 32086 && 
b[32087] == 32087 && 
b[32088] == 32088 && 
b[32089] == 32089 && 
b[32090] == 32090 && 
b[32091] == 32091 && 
b[32092] == 32092 && 
b[32093] == 32093 && 
b[32094] == 32094 && 
b[32095] == 32095 && 
b[32096] == 32096 && 
b[32097] == 32097 && 
b[32098] == 32098 && 
b[32099] == 32099 && 
b[32100] == 32100 && 
b[32101] == 32101 && 
b[32102] == 32102 && 
b[32103] == 32103 && 
b[32104] == 32104 && 
b[32105] == 32105 && 
b[32106] == 32106 && 
b[32107] == 32107 && 
b[32108] == 32108 && 
b[32109] == 32109 && 
b[32110] == 32110 && 
b[32111] == 32111 && 
b[32112] == 32112 && 
b[32113] == 32113 && 
b[32114] == 32114 && 
b[32115] == 32115 && 
b[32116] == 32116 && 
b[32117] == 32117 && 
b[32118] == 32118 && 
b[32119] == 32119 && 
b[32120] == 32120 && 
b[32121] == 32121 && 
b[32122] == 32122 && 
b[32123] == 32123 && 
b[32124] == 32124 && 
b[32125] == 32125 && 
b[32126] == 32126 && 
b[32127] == 32127 && 
b[32128] == 32128 && 
b[32129] == 32129 && 
b[32130] == 32130 && 
b[32131] == 32131 && 
b[32132] == 32132 && 
b[32133] == 32133 && 
b[32134] == 32134 && 
b[32135] == 32135 && 
b[32136] == 32136 && 
b[32137] == 32137 && 
b[32138] == 32138 && 
b[32139] == 32139 && 
b[32140] == 32140 && 
b[32141] == 32141 && 
b[32142] == 32142 && 
b[32143] == 32143 && 
b[32144] == 32144 && 
b[32145] == 32145 && 
b[32146] == 32146 && 
b[32147] == 32147 && 
b[32148] == 32148 && 
b[32149] == 32149 && 
b[32150] == 32150 && 
b[32151] == 32151 && 
b[32152] == 32152 && 
b[32153] == 32153 && 
b[32154] == 32154 && 
b[32155] == 32155 && 
b[32156] == 32156 && 
b[32157] == 32157 && 
b[32158] == 32158 && 
b[32159] == 32159 && 
b[32160] == 32160 && 
b[32161] == 32161 && 
b[32162] == 32162 && 
b[32163] == 32163 && 
b[32164] == 32164 && 
b[32165] == 32165 && 
b[32166] == 32166 && 
b[32167] == 32167 && 
b[32168] == 32168 && 
b[32169] == 32169 && 
b[32170] == 32170 && 
b[32171] == 32171 && 
b[32172] == 32172 && 
b[32173] == 32173 && 
b[32174] == 32174 && 
b[32175] == 32175 && 
b[32176] == 32176 && 
b[32177] == 32177 && 
b[32178] == 32178 && 
b[32179] == 32179 && 
b[32180] == 32180 && 
b[32181] == 32181 && 
b[32182] == 32182 && 
b[32183] == 32183 && 
b[32184] == 32184 && 
b[32185] == 32185 && 
b[32186] == 32186 && 
b[32187] == 32187 && 
b[32188] == 32188 && 
b[32189] == 32189 && 
b[32190] == 32190 && 
b[32191] == 32191 && 
b[32192] == 32192 && 
b[32193] == 32193 && 
b[32194] == 32194 && 
b[32195] == 32195 && 
b[32196] == 32196 && 
b[32197] == 32197 && 
b[32198] == 32198 && 
b[32199] == 32199 && 
b[32200] == 32200 && 
b[32201] == 32201 && 
b[32202] == 32202 && 
b[32203] == 32203 && 
b[32204] == 32204 && 
b[32205] == 32205 && 
b[32206] == 32206 && 
b[32207] == 32207 && 
b[32208] == 32208 && 
b[32209] == 32209 && 
b[32210] == 32210 && 
b[32211] == 32211 && 
b[32212] == 32212 && 
b[32213] == 32213 && 
b[32214] == 32214 && 
b[32215] == 32215 && 
b[32216] == 32216 && 
b[32217] == 32217 && 
b[32218] == 32218 && 
b[32219] == 32219 && 
b[32220] == 32220 && 
b[32221] == 32221 && 
b[32222] == 32222 && 
b[32223] == 32223 && 
b[32224] == 32224 && 
b[32225] == 32225 && 
b[32226] == 32226 && 
b[32227] == 32227 && 
b[32228] == 32228 && 
b[32229] == 32229 && 
b[32230] == 32230 && 
b[32231] == 32231 && 
b[32232] == 32232 && 
b[32233] == 32233 && 
b[32234] == 32234 && 
b[32235] == 32235 && 
b[32236] == 32236 && 
b[32237] == 32237 && 
b[32238] == 32238 && 
b[32239] == 32239 && 
b[32240] == 32240 && 
b[32241] == 32241 && 
b[32242] == 32242 && 
b[32243] == 32243 && 
b[32244] == 32244 && 
b[32245] == 32245 && 
b[32246] == 32246 && 
b[32247] == 32247 && 
b[32248] == 32248 && 
b[32249] == 32249 && 
b[32250] == 32250 && 
b[32251] == 32251 && 
b[32252] == 32252 && 
b[32253] == 32253 && 
b[32254] == 32254 && 
b[32255] == 32255 && 
b[32256] == 32256 && 
b[32257] == 32257 && 
b[32258] == 32258 && 
b[32259] == 32259 && 
b[32260] == 32260 && 
b[32261] == 32261 && 
b[32262] == 32262 && 
b[32263] == 32263 && 
b[32264] == 32264 && 
b[32265] == 32265 && 
b[32266] == 32266 && 
b[32267] == 32267 && 
b[32268] == 32268 && 
b[32269] == 32269 && 
b[32270] == 32270 && 
b[32271] == 32271 && 
b[32272] == 32272 && 
b[32273] == 32273 && 
b[32274] == 32274 && 
b[32275] == 32275 && 
b[32276] == 32276 && 
b[32277] == 32277 && 
b[32278] == 32278 && 
b[32279] == 32279 && 
b[32280] == 32280 && 
b[32281] == 32281 && 
b[32282] == 32282 && 
b[32283] == 32283 && 
b[32284] == 32284 && 
b[32285] == 32285 && 
b[32286] == 32286 && 
b[32287] == 32287 && 
b[32288] == 32288 && 
b[32289] == 32289 && 
b[32290] == 32290 && 
b[32291] == 32291 && 
b[32292] == 32292 && 
b[32293] == 32293 && 
b[32294] == 32294 && 
b[32295] == 32295 && 
b[32296] == 32296 && 
b[32297] == 32297 && 
b[32298] == 32298 && 
b[32299] == 32299 && 
b[32300] == 32300 && 
b[32301] == 32301 && 
b[32302] == 32302 && 
b[32303] == 32303 && 
b[32304] == 32304 && 
b[32305] == 32305 && 
b[32306] == 32306 && 
b[32307] == 32307 && 
b[32308] == 32308 && 
b[32309] == 32309 && 
b[32310] == 32310 && 
b[32311] == 32311 && 
b[32312] == 32312 && 
b[32313] == 32313 && 
b[32314] == 32314 && 
b[32315] == 32315 && 
b[32316] == 32316 && 
b[32317] == 32317 && 
b[32318] == 32318 && 
b[32319] == 32319 && 
b[32320] == 32320 && 
b[32321] == 32321 && 
b[32322] == 32322 && 
b[32323] == 32323 && 
b[32324] == 32324 && 
b[32325] == 32325 && 
b[32326] == 32326 && 
b[32327] == 32327 && 
b[32328] == 32328 && 
b[32329] == 32329 && 
b[32330] == 32330 && 
b[32331] == 32331 && 
b[32332] == 32332 && 
b[32333] == 32333 && 
b[32334] == 32334 && 
b[32335] == 32335 && 
b[32336] == 32336 && 
b[32337] == 32337 && 
b[32338] == 32338 && 
b[32339] == 32339 && 
b[32340] == 32340 && 
b[32341] == 32341 && 
b[32342] == 32342 && 
b[32343] == 32343 && 
b[32344] == 32344 && 
b[32345] == 32345 && 
b[32346] == 32346 && 
b[32347] == 32347 && 
b[32348] == 32348 && 
b[32349] == 32349 && 
b[32350] == 32350 && 
b[32351] == 32351 && 
b[32352] == 32352 && 
b[32353] == 32353 && 
b[32354] == 32354 && 
b[32355] == 32355 && 
b[32356] == 32356 && 
b[32357] == 32357 && 
b[32358] == 32358 && 
b[32359] == 32359 && 
b[32360] == 32360 && 
b[32361] == 32361 && 
b[32362] == 32362 && 
b[32363] == 32363 && 
b[32364] == 32364 && 
b[32365] == 32365 && 
b[32366] == 32366 && 
b[32367] == 32367 && 
b[32368] == 32368 && 
b[32369] == 32369 && 
b[32370] == 32370 && 
b[32371] == 32371 && 
b[32372] == 32372 && 
b[32373] == 32373 && 
b[32374] == 32374 && 
b[32375] == 32375 && 
b[32376] == 32376 && 
b[32377] == 32377 && 
b[32378] == 32378 && 
b[32379] == 32379 && 
b[32380] == 32380 && 
b[32381] == 32381 && 
b[32382] == 32382 && 
b[32383] == 32383 && 
b[32384] == 32384 && 
b[32385] == 32385 && 
b[32386] == 32386 && 
b[32387] == 32387 && 
b[32388] == 32388 && 
b[32389] == 32389 && 
b[32390] == 32390 && 
b[32391] == 32391 && 
b[32392] == 32392 && 
b[32393] == 32393 && 
b[32394] == 32394 && 
b[32395] == 32395 && 
b[32396] == 32396 && 
b[32397] == 32397 && 
b[32398] == 32398 && 
b[32399] == 32399 && 
b[32400] == 32400 && 
b[32401] == 32401 && 
b[32402] == 32402 && 
b[32403] == 32403 && 
b[32404] == 32404 && 
b[32405] == 32405 && 
b[32406] == 32406 && 
b[32407] == 32407 && 
b[32408] == 32408 && 
b[32409] == 32409 && 
b[32410] == 32410 && 
b[32411] == 32411 && 
b[32412] == 32412 && 
b[32413] == 32413 && 
b[32414] == 32414 && 
b[32415] == 32415 && 
b[32416] == 32416 && 
b[32417] == 32417 && 
b[32418] == 32418 && 
b[32419] == 32419 && 
b[32420] == 32420 && 
b[32421] == 32421 && 
b[32422] == 32422 && 
b[32423] == 32423 && 
b[32424] == 32424 && 
b[32425] == 32425 && 
b[32426] == 32426 && 
b[32427] == 32427 && 
b[32428] == 32428 && 
b[32429] == 32429 && 
b[32430] == 32430 && 
b[32431] == 32431 && 
b[32432] == 32432 && 
b[32433] == 32433 && 
b[32434] == 32434 && 
b[32435] == 32435 && 
b[32436] == 32436 && 
b[32437] == 32437 && 
b[32438] == 32438 && 
b[32439] == 32439 && 
b[32440] == 32440 && 
b[32441] == 32441 && 
b[32442] == 32442 && 
b[32443] == 32443 && 
b[32444] == 32444 && 
b[32445] == 32445 && 
b[32446] == 32446 && 
b[32447] == 32447 && 
b[32448] == 32448 && 
b[32449] == 32449 && 
b[32450] == 32450 && 
b[32451] == 32451 && 
b[32452] == 32452 && 
b[32453] == 32453 && 
b[32454] == 32454 && 
b[32455] == 32455 && 
b[32456] == 32456 && 
b[32457] == 32457 && 
b[32458] == 32458 && 
b[32459] == 32459 && 
b[32460] == 32460 && 
b[32461] == 32461 && 
b[32462] == 32462 && 
b[32463] == 32463 && 
b[32464] == 32464 && 
b[32465] == 32465 && 
b[32466] == 32466 && 
b[32467] == 32467 && 
b[32468] == 32468 && 
b[32469] == 32469 && 
b[32470] == 32470 && 
b[32471] == 32471 && 
b[32472] == 32472 && 
b[32473] == 32473 && 
b[32474] == 32474 && 
b[32475] == 32475 && 
b[32476] == 32476 && 
b[32477] == 32477 && 
b[32478] == 32478 && 
b[32479] == 32479 && 
b[32480] == 32480 && 
b[32481] == 32481 && 
b[32482] == 32482 && 
b[32483] == 32483 && 
b[32484] == 32484 && 
b[32485] == 32485 && 
b[32486] == 32486 && 
b[32487] == 32487 && 
b[32488] == 32488 && 
b[32489] == 32489 && 
b[32490] == 32490 && 
b[32491] == 32491 && 
b[32492] == 32492 && 
b[32493] == 32493 && 
b[32494] == 32494 && 
b[32495] == 32495 && 
b[32496] == 32496 && 
b[32497] == 32497 && 
b[32498] == 32498 && 
b[32499] == 32499 && 
b[32500] == 32500 && 
b[32501] == 32501 && 
b[32502] == 32502 && 
b[32503] == 32503 && 
b[32504] == 32504 && 
b[32505] == 32505 && 
b[32506] == 32506 && 
b[32507] == 32507 && 
b[32508] == 32508 && 
b[32509] == 32509 && 
b[32510] == 32510 && 
b[32511] == 32511 && 
b[32512] == 32512 && 
b[32513] == 32513 && 
b[32514] == 32514 && 
b[32515] == 32515 && 
b[32516] == 32516 && 
b[32517] == 32517 && 
b[32518] == 32518 && 
b[32519] == 32519 && 
b[32520] == 32520 && 
b[32521] == 32521 && 
b[32522] == 32522 && 
b[32523] == 32523 && 
b[32524] == 32524 && 
b[32525] == 32525 && 
b[32526] == 32526 && 
b[32527] == 32527 && 
b[32528] == 32528 && 
b[32529] == 32529 && 
b[32530] == 32530 && 
b[32531] == 32531 && 
b[32532] == 32532 && 
b[32533] == 32533 && 
b[32534] == 32534 && 
b[32535] == 32535 && 
b[32536] == 32536 && 
b[32537] == 32537 && 
b[32538] == 32538 && 
b[32539] == 32539 && 
b[32540] == 32540 && 
b[32541] == 32541 && 
b[32542] == 32542 && 
b[32543] == 32543 && 
b[32544] == 32544 && 
b[32545] == 32545 && 
b[32546] == 32546 && 
b[32547] == 32547 && 
b[32548] == 32548 && 
b[32549] == 32549 && 
b[32550] == 32550 && 
b[32551] == 32551 && 
b[32552] == 32552 && 
b[32553] == 32553 && 
b[32554] == 32554 && 
b[32555] == 32555 && 
b[32556] == 32556 && 
b[32557] == 32557 && 
b[32558] == 32558 && 
b[32559] == 32559 && 
b[32560] == 32560 && 
b[32561] == 32561 && 
b[32562] == 32562 && 
b[32563] == 32563 && 
b[32564] == 32564 && 
b[32565] == 32565 && 
b[32566] == 32566 && 
b[32567] == 32567 && 
b[32568] == 32568 && 
b[32569] == 32569 && 
b[32570] == 32570 && 
b[32571] == 32571 && 
b[32572] == 32572 && 
b[32573] == 32573 && 
b[32574] == 32574 && 
b[32575] == 32575 && 
b[32576] == 32576 && 
b[32577] == 32577 && 
b[32578] == 32578 && 
b[32579] == 32579 && 
b[32580] == 32580 && 
b[32581] == 32581 && 
b[32582] == 32582 && 
b[32583] == 32583 && 
b[32584] == 32584 && 
b[32585] == 32585 && 
b[32586] == 32586 && 
b[32587] == 32587 && 
b[32588] == 32588 && 
b[32589] == 32589 && 
b[32590] == 32590 && 
b[32591] == 32591 && 
b[32592] == 32592 && 
b[32593] == 32593 && 
b[32594] == 32594 && 
b[32595] == 32595 && 
b[32596] == 32596 && 
b[32597] == 32597 && 
b[32598] == 32598 && 
b[32599] == 32599 && 
b[32600] == 32600 && 
b[32601] == 32601 && 
b[32602] == 32602 && 
b[32603] == 32603 && 
b[32604] == 32604 && 
b[32605] == 32605 && 
b[32606] == 32606 && 
b[32607] == 32607 && 
b[32608] == 32608 && 
b[32609] == 32609 && 
b[32610] == 32610 && 
b[32611] == 32611 && 
b[32612] == 32612 && 
b[32613] == 32613 && 
b[32614] == 32614 && 
b[32615] == 32615 && 
b[32616] == 32616 && 
b[32617] == 32617 && 
b[32618] == 32618 && 
b[32619] == 32619 && 
b[32620] == 32620 && 
b[32621] == 32621 && 
b[32622] == 32622 && 
b[32623] == 32623 && 
b[32624] == 32624 && 
b[32625] == 32625 && 
b[32626] == 32626 && 
b[32627] == 32627 && 
b[32628] == 32628 && 
b[32629] == 32629 && 
b[32630] == 32630 && 
b[32631] == 32631 && 
b[32632] == 32632 && 
b[32633] == 32633 && 
b[32634] == 32634 && 
b[32635] == 32635 && 
b[32636] == 32636 && 
b[32637] == 32637 && 
b[32638] == 32638 && 
b[32639] == 32639 && 
b[32640] == 32640 && 
b[32641] == 32641 && 
b[32642] == 32642 && 
b[32643] == 32643 && 
b[32644] == 32644 && 
b[32645] == 32645 && 
b[32646] == 32646 && 
b[32647] == 32647 && 
b[32648] == 32648 && 
b[32649] == 32649 && 
b[32650] == 32650 && 
b[32651] == 32651 && 
b[32652] == 32652 && 
b[32653] == 32653 && 
b[32654] == 32654 && 
b[32655] == 32655 && 
b[32656] == 32656 && 
b[32657] == 32657 && 
b[32658] == 32658 && 
b[32659] == 32659 && 
b[32660] == 32660 && 
b[32661] == 32661 && 
b[32662] == 32662 && 
b[32663] == 32663 && 
b[32664] == 32664 && 
b[32665] == 32665 && 
b[32666] == 32666 && 
b[32667] == 32667 && 
b[32668] == 32668 && 
b[32669] == 32669 && 
b[32670] == 32670 && 
b[32671] == 32671 && 
b[32672] == 32672 && 
b[32673] == 32673 && 
b[32674] == 32674 && 
b[32675] == 32675 && 
b[32676] == 32676 && 
b[32677] == 32677 && 
b[32678] == 32678 && 
b[32679] == 32679 && 
b[32680] == 32680 && 
b[32681] == 32681 && 
b[32682] == 32682 && 
b[32683] == 32683 && 
b[32684] == 32684 && 
b[32685] == 32685 && 
b[32686] == 32686 && 
b[32687] == 32687 && 
b[32688] == 32688 && 
b[32689] == 32689 && 
b[32690] == 32690 && 
b[32691] == 32691 && 
b[32692] == 32692 && 
b[32693] == 32693 && 
b[32694] == 32694 && 
b[32695] == 32695 && 
b[32696] == 32696 && 
b[32697] == 32697 && 
b[32698] == 32698 && 
b[32699] == 32699 && 
b[32700] == 32700 && 
b[32701] == 32701 && 
b[32702] == 32702 && 
b[32703] == 32703 && 
b[32704] == 32704 && 
b[32705] == 32705 && 
b[32706] == 32706 && 
b[32707] == 32707 && 
b[32708] == 32708 && 
b[32709] == 32709 && 
b[32710] == 32710 && 
b[32711] == 32711 && 
b[32712] == 32712 && 
b[32713] == 32713 && 
b[32714] == 32714 && 
b[32715] == 32715 && 
b[32716] == 32716 && 
b[32717] == 32717 && 
b[32718] == 32718 && 
b[32719] == 32719 && 
b[32720] == 32720 && 
b[32721] == 32721 && 
b[32722] == 32722 && 
b[32723] == 32723 && 
b[32724] == 32724 && 
b[32725] == 32725 && 
b[32726] == 32726 && 
b[32727] == 32727 && 
b[32728] == 32728 && 
b[32729] == 32729 && 
b[32730] == 32730 && 
b[32731] == 32731 && 
b[32732] == 32732 && 
b[32733] == 32733 && 
b[32734] == 32734 && 
b[32735] == 32735 && 
b[32736] == 32736 && 
b[32737] == 32737 && 
b[32738] == 32738 && 
b[32739] == 32739 && 
b[32740] == 32740 && 
b[32741] == 32741 && 
b[32742] == 32742 && 
b[32743] == 32743 && 
b[32744] == 32744 && 
b[32745] == 32745 && 
b[32746] == 32746 && 
b[32747] == 32747 && 
b[32748] == 32748 && 
b[32749] == 32749 && 
b[32750] == 32750 && 
b[32751] == 32751 && 
b[32752] == 32752 && 
b[32753] == 32753 && 
b[32754] == 32754 && 
b[32755] == 32755 && 
b[32756] == 32756 && 
b[32757] == 32757 && 
b[32758] == 32758 && 
b[32759] == 32759 && 
b[32760] == 32760 && 
b[32761] == 32761 && 
b[32762] == 32762 && 
b[32763] == 32763 && 
b[32764] == 32764 && 
b[32765] == 32765 && 
b[32766] == 32766 && 
b[32767] == 32767 && 
b[32768] == 32768 && 
b[32769] == 32769 && 
b[32770] == 32770 && 
b[32771] == 32771 && 
b[32772] == 32772 && 
b[32773] == 32773 && 
b[32774] == 32774 && 
b[32775] == 32775 && 
b[32776] == 32776 && 
b[32777] == 32777 && 
b[32778] == 32778 && 
b[32779] == 32779 && 
b[32780] == 32780 && 
b[32781] == 32781 && 
b[32782] == 32782 && 
b[32783] == 32783 && 
b[32784] == 32784 && 
b[32785] == 32785 && 
b[32786] == 32786 && 
b[32787] == 32787 && 
b[32788] == 32788 && 
b[32789] == 32789 && 
b[32790] == 32790 && 
b[32791] == 32791 && 
b[32792] == 32792 && 
b[32793] == 32793 && 
b[32794] == 32794 && 
b[32795] == 32795 && 
b[32796] == 32796 && 
b[32797] == 32797 && 
b[32798] == 32798 && 
b[32799] == 32799 && 
b[32800] == 32800 && 
b[32801] == 32801 && 
b[32802] == 32802 && 
b[32803] == 32803 && 
b[32804] == 32804 && 
b[32805] == 32805 && 
b[32806] == 32806 && 
b[32807] == 32807 && 
b[32808] == 32808 && 
b[32809] == 32809 && 
b[32810] == 32810 && 
b[32811] == 32811 && 
b[32812] == 32812 && 
b[32813] == 32813 && 
b[32814] == 32814 && 
b[32815] == 32815 && 
b[32816] == 32816 && 
b[32817] == 32817 && 
b[32818] == 32818 && 
b[32819] == 32819 && 
b[32820] == 32820 && 
b[32821] == 32821 && 
b[32822] == 32822 && 
b[32823] == 32823 && 
b[32824] == 32824 && 
b[32825] == 32825 && 
b[32826] == 32826 && 
b[32827] == 32827 && 
b[32828] == 32828 && 
b[32829] == 32829 && 
b[32830] == 32830 && 
b[32831] == 32831 && 
b[32832] == 32832 && 
b[32833] == 32833 && 
b[32834] == 32834 && 
b[32835] == 32835 && 
b[32836] == 32836 && 
b[32837] == 32837 && 
b[32838] == 32838 && 
b[32839] == 32839 && 
b[32840] == 32840 && 
b[32841] == 32841 && 
b[32842] == 32842 && 
b[32843] == 32843 && 
b[32844] == 32844 && 
b[32845] == 32845 && 
b[32846] == 32846 && 
b[32847] == 32847 && 
b[32848] == 32848 && 
b[32849] == 32849 && 
b[32850] == 32850 && 
b[32851] == 32851 && 
b[32852] == 32852 && 
b[32853] == 32853 && 
b[32854] == 32854 && 
b[32855] == 32855 && 
b[32856] == 32856 && 
b[32857] == 32857 && 
b[32858] == 32858 && 
b[32859] == 32859 && 
b[32860] == 32860 && 
b[32861] == 32861 && 
b[32862] == 32862 && 
b[32863] == 32863 && 
b[32864] == 32864 && 
b[32865] == 32865 && 
b[32866] == 32866 && 
b[32867] == 32867 && 
b[32868] == 32868 && 
b[32869] == 32869 && 
b[32870] == 32870 && 
b[32871] == 32871 && 
b[32872] == 32872 && 
b[32873] == 32873 && 
b[32874] == 32874 && 
b[32875] == 32875 && 
b[32876] == 32876 && 
b[32877] == 32877 && 
b[32878] == 32878 && 
b[32879] == 32879 && 
b[32880] == 32880 && 
b[32881] == 32881 && 
b[32882] == 32882 && 
b[32883] == 32883 && 
b[32884] == 32884 && 
b[32885] == 32885 && 
b[32886] == 32886 && 
b[32887] == 32887 && 
b[32888] == 32888 && 
b[32889] == 32889 && 
b[32890] == 32890 && 
b[32891] == 32891 && 
b[32892] == 32892 && 
b[32893] == 32893 && 
b[32894] == 32894 && 
b[32895] == 32895 && 
b[32896] == 32896 && 
b[32897] == 32897 && 
b[32898] == 32898 && 
b[32899] == 32899 && 
b[32900] == 32900 && 
b[32901] == 32901 && 
b[32902] == 32902 && 
b[32903] == 32903 && 
b[32904] == 32904 && 
b[32905] == 32905 && 
b[32906] == 32906 && 
b[32907] == 32907 && 
b[32908] == 32908 && 
b[32909] == 32909 && 
b[32910] == 32910 && 
b[32911] == 32911 && 
b[32912] == 32912 && 
b[32913] == 32913 && 
b[32914] == 32914 && 
b[32915] == 32915 && 
b[32916] == 32916 && 
b[32917] == 32917 && 
b[32918] == 32918 && 
b[32919] == 32919 && 
b[32920] == 32920 && 
b[32921] == 32921 && 
b[32922] == 32922 && 
b[32923] == 32923 && 
b[32924] == 32924 && 
b[32925] == 32925 && 
b[32926] == 32926 && 
b[32927] == 32927 && 
b[32928] == 32928 && 
b[32929] == 32929 && 
b[32930] == 32930 && 
b[32931] == 32931 && 
b[32932] == 32932 && 
b[32933] == 32933 && 
b[32934] == 32934 && 
b[32935] == 32935 && 
b[32936] == 32936 && 
b[32937] == 32937 && 
b[32938] == 32938 && 
b[32939] == 32939 && 
b[32940] == 32940 && 
b[32941] == 32941 && 
b[32942] == 32942 && 
b[32943] == 32943 && 
b[32944] == 32944 && 
b[32945] == 32945 && 
b[32946] == 32946 && 
b[32947] == 32947 && 
b[32948] == 32948 && 
b[32949] == 32949 && 
b[32950] == 32950 && 
b[32951] == 32951 && 
b[32952] == 32952 && 
b[32953] == 32953 && 
b[32954] == 32954 && 
b[32955] == 32955 && 
b[32956] == 32956 && 
b[32957] == 32957 && 
b[32958] == 32958 && 
b[32959] == 32959 && 
b[32960] == 32960 && 
b[32961] == 32961 && 
b[32962] == 32962 && 
b[32963] == 32963 && 
b[32964] == 32964 && 
b[32965] == 32965 && 
b[32966] == 32966 && 
b[32967] == 32967 && 
b[32968] == 32968 && 
b[32969] == 32969 && 
b[32970] == 32970 && 
b[32971] == 32971 && 
b[32972] == 32972 && 
b[32973] == 32973 && 
b[32974] == 32974 && 
b[32975] == 32975 && 
b[32976] == 32976 && 
b[32977] == 32977 && 
b[32978] == 32978 && 
b[32979] == 32979 && 
b[32980] == 32980 && 
b[32981] == 32981 && 
b[32982] == 32982 && 
b[32983] == 32983 && 
b[32984] == 32984 && 
b[32985] == 32985 && 
b[32986] == 32986 && 
b[32987] == 32987 && 
b[32988] == 32988 && 
b[32989] == 32989 && 
b[32990] == 32990 && 
b[32991] == 32991 && 
b[32992] == 32992 && 
b[32993] == 32993 && 
b[32994] == 32994 && 
b[32995] == 32995 && 
b[32996] == 32996 && 
b[32997] == 32997 && 
b[32998] == 32998 && 
b[32999] == 32999 && 
b[33000] == 33000 && 
b[33001] == 33001 && 
b[33002] == 33002 && 
b[33003] == 33003 && 
b[33004] == 33004 && 
b[33005] == 33005 && 
b[33006] == 33006 && 
b[33007] == 33007 && 
b[33008] == 33008 && 
b[33009] == 33009 && 
b[33010] == 33010 && 
b[33011] == 33011 && 
b[33012] == 33012 && 
b[33013] == 33013 && 
b[33014] == 33014 && 
b[33015] == 33015 && 
b[33016] == 33016 && 
b[33017] == 33017 && 
b[33018] == 33018 && 
b[33019] == 33019 && 
b[33020] == 33020 && 
b[33021] == 33021 && 
b[33022] == 33022 && 
b[33023] == 33023 && 
b[33024] == 33024 && 
b[33025] == 33025 && 
b[33026] == 33026 && 
b[33027] == 33027 && 
b[33028] == 33028 && 
b[33029] == 33029 && 
b[33030] == 33030 && 
b[33031] == 33031 && 
b[33032] == 33032 && 
b[33033] == 33033 && 
b[33034] == 33034 && 
b[33035] == 33035 && 
b[33036] == 33036 && 
b[33037] == 33037 && 
b[33038] == 33038 && 
b[33039] == 33039 && 
b[33040] == 33040 && 
b[33041] == 33041 && 
b[33042] == 33042 && 
b[33043] == 33043 && 
b[33044] == 33044 && 
b[33045] == 33045 && 
b[33046] == 33046 && 
b[33047] == 33047 && 
b[33048] == 33048 && 
b[33049] == 33049 && 
b[33050] == 33050 && 
b[33051] == 33051 && 
b[33052] == 33052 && 
b[33053] == 33053 && 
b[33054] == 33054 && 
b[33055] == 33055 && 
b[33056] == 33056 && 
b[33057] == 33057 && 
b[33058] == 33058 && 
b[33059] == 33059 && 
b[33060] == 33060 && 
b[33061] == 33061 && 
b[33062] == 33062 && 
b[33063] == 33063 && 
b[33064] == 33064 && 
b[33065] == 33065 && 
b[33066] == 33066 && 
b[33067] == 33067 && 
b[33068] == 33068 && 
b[33069] == 33069 && 
b[33070] == 33070 && 
b[33071] == 33071 && 
b[33072] == 33072 && 
b[33073] == 33073 && 
b[33074] == 33074 && 
b[33075] == 33075 && 
b[33076] == 33076 && 
b[33077] == 33077 && 
b[33078] == 33078 && 
b[33079] == 33079 && 
b[33080] == 33080 && 
b[33081] == 33081 && 
b[33082] == 33082 && 
b[33083] == 33083 && 
b[33084] == 33084 && 
b[33085] == 33085 && 
b[33086] == 33086 && 
b[33087] == 33087 && 
b[33088] == 33088 && 
b[33089] == 33089 && 
b[33090] == 33090 && 
b[33091] == 33091 && 
b[33092] == 33092 && 
b[33093] == 33093 && 
b[33094] == 33094 && 
b[33095] == 33095 && 
b[33096] == 33096 && 
b[33097] == 33097 && 
b[33098] == 33098 && 
b[33099] == 33099 && 
b[33100] == 33100 && 
b[33101] == 33101 && 
b[33102] == 33102 && 
b[33103] == 33103 && 
b[33104] == 33104 && 
b[33105] == 33105 && 
b[33106] == 33106 && 
b[33107] == 33107 && 
b[33108] == 33108 && 
b[33109] == 33109 && 
b[33110] == 33110 && 
b[33111] == 33111 && 
b[33112] == 33112 && 
b[33113] == 33113 && 
b[33114] == 33114 && 
b[33115] == 33115 && 
b[33116] == 33116 && 
b[33117] == 33117 && 
b[33118] == 33118 && 
b[33119] == 33119 && 
b[33120] == 33120 && 
b[33121] == 33121 && 
b[33122] == 33122 && 
b[33123] == 33123 && 
b[33124] == 33124 && 
b[33125] == 33125 && 
b[33126] == 33126 && 
b[33127] == 33127 && 
b[33128] == 33128 && 
b[33129] == 33129 && 
b[33130] == 33130 && 
b[33131] == 33131 && 
b[33132] == 33132 && 
b[33133] == 33133 && 
b[33134] == 33134 && 
b[33135] == 33135 && 
b[33136] == 33136 && 
b[33137] == 33137 && 
b[33138] == 33138 && 
b[33139] == 33139 && 
b[33140] == 33140 && 
b[33141] == 33141 && 
b[33142] == 33142 && 
b[33143] == 33143 && 
b[33144] == 33144 && 
b[33145] == 33145 && 
b[33146] == 33146 && 
b[33147] == 33147 && 
b[33148] == 33148 && 
b[33149] == 33149 && 
b[33150] == 33150 && 
b[33151] == 33151 && 
b[33152] == 33152 && 
b[33153] == 33153 && 
b[33154] == 33154 && 
b[33155] == 33155 && 
b[33156] == 33156 && 
b[33157] == 33157 && 
b[33158] == 33158 && 
b[33159] == 33159 && 
b[33160] == 33160 && 
b[33161] == 33161 && 
b[33162] == 33162 && 
b[33163] == 33163 && 
b[33164] == 33164 && 
b[33165] == 33165 && 
b[33166] == 33166 && 
b[33167] == 33167 && 
b[33168] == 33168 && 
b[33169] == 33169 && 
b[33170] == 33170 && 
b[33171] == 33171 && 
b[33172] == 33172 && 
b[33173] == 33173 && 
b[33174] == 33174 && 
b[33175] == 33175 && 
b[33176] == 33176 && 
b[33177] == 33177 && 
b[33178] == 33178 && 
b[33179] == 33179 && 
b[33180] == 33180 && 
b[33181] == 33181 && 
b[33182] == 33182 && 
b[33183] == 33183 && 
b[33184] == 33184 && 
b[33185] == 33185 && 
b[33186] == 33186 && 
b[33187] == 33187 && 
b[33188] == 33188 && 
b[33189] == 33189 && 
b[33190] == 33190 && 
b[33191] == 33191 && 
b[33192] == 33192 && 
b[33193] == 33193 && 
b[33194] == 33194 && 
b[33195] == 33195 && 
b[33196] == 33196 && 
b[33197] == 33197 && 
b[33198] == 33198 && 
b[33199] == 33199 && 
b[33200] == 33200 && 
b[33201] == 33201 && 
b[33202] == 33202 && 
b[33203] == 33203 && 
b[33204] == 33204 && 
b[33205] == 33205 && 
b[33206] == 33206 && 
b[33207] == 33207 && 
b[33208] == 33208 && 
b[33209] == 33209 && 
b[33210] == 33210 && 
b[33211] == 33211 && 
b[33212] == 33212 && 
b[33213] == 33213 && 
b[33214] == 33214 && 
b[33215] == 33215 && 
b[33216] == 33216 && 
b[33217] == 33217 && 
b[33218] == 33218 && 
b[33219] == 33219 && 
b[33220] == 33220 && 
b[33221] == 33221 && 
b[33222] == 33222 && 
b[33223] == 33223 && 
b[33224] == 33224 && 
b[33225] == 33225 && 
b[33226] == 33226 && 
b[33227] == 33227 && 
b[33228] == 33228 && 
b[33229] == 33229 && 
b[33230] == 33230 && 
b[33231] == 33231 && 
b[33232] == 33232 && 
b[33233] == 33233 && 
b[33234] == 33234 && 
b[33235] == 33235 && 
b[33236] == 33236 && 
b[33237] == 33237 && 
b[33238] == 33238 && 
b[33239] == 33239 && 
b[33240] == 33240 && 
b[33241] == 33241 && 
b[33242] == 33242 && 
b[33243] == 33243 && 
b[33244] == 33244 && 
b[33245] == 33245 && 
b[33246] == 33246 && 
b[33247] == 33247 && 
b[33248] == 33248 && 
b[33249] == 33249 && 
b[33250] == 33250 && 
b[33251] == 33251 && 
b[33252] == 33252 && 
b[33253] == 33253 && 
b[33254] == 33254 && 
b[33255] == 33255 && 
b[33256] == 33256 && 
b[33257] == 33257 && 
b[33258] == 33258 && 
b[33259] == 33259 && 
b[33260] == 33260 && 
b[33261] == 33261 && 
b[33262] == 33262 && 
b[33263] == 33263 && 
b[33264] == 33264 && 
b[33265] == 33265 && 
b[33266] == 33266 && 
b[33267] == 33267 && 
b[33268] == 33268 && 
b[33269] == 33269 && 
b[33270] == 33270 && 
b[33271] == 33271 && 
b[33272] == 33272 && 
b[33273] == 33273 && 
b[33274] == 33274 && 
b[33275] == 33275 && 
b[33276] == 33276 && 
b[33277] == 33277 && 
b[33278] == 33278 && 
b[33279] == 33279 && 
b[33280] == 33280 && 
b[33281] == 33281 && 
b[33282] == 33282 && 
b[33283] == 33283 && 
b[33284] == 33284 && 
b[33285] == 33285 && 
b[33286] == 33286 && 
b[33287] == 33287 && 
b[33288] == 33288 && 
b[33289] == 33289 && 
b[33290] == 33290 && 
b[33291] == 33291 && 
b[33292] == 33292 && 
b[33293] == 33293 && 
b[33294] == 33294 && 
b[33295] == 33295 && 
b[33296] == 33296 && 
b[33297] == 33297 && 
b[33298] == 33298 && 
b[33299] == 33299 && 
b[33300] == 33300 && 
b[33301] == 33301 && 
b[33302] == 33302 && 
b[33303] == 33303 && 
b[33304] == 33304 && 
b[33305] == 33305 && 
b[33306] == 33306 && 
b[33307] == 33307 && 
b[33308] == 33308 && 
b[33309] == 33309 && 
b[33310] == 33310 && 
b[33311] == 33311 && 
b[33312] == 33312 && 
b[33313] == 33313 && 
b[33314] == 33314 && 
b[33315] == 33315 && 
b[33316] == 33316 && 
b[33317] == 33317 && 
b[33318] == 33318 && 
b[33319] == 33319 && 
b[33320] == 33320 && 
b[33321] == 33321 && 
b[33322] == 33322 && 
b[33323] == 33323 && 
b[33324] == 33324 && 
b[33325] == 33325 && 
b[33326] == 33326 && 
b[33327] == 33327 && 
b[33328] == 33328 && 
b[33329] == 33329 && 
b[33330] == 33330 && 
b[33331] == 33331 && 
b[33332] == 33332 && 
b[33333] == 33333 && 
b[33334] == 33334 && 
b[33335] == 33335 && 
b[33336] == 33336 && 
b[33337] == 33337 && 
b[33338] == 33338 && 
b[33339] == 33339 && 
b[33340] == 33340 && 
b[33341] == 33341 && 
b[33342] == 33342 && 
b[33343] == 33343 && 
b[33344] == 33344 && 
b[33345] == 33345 && 
b[33346] == 33346 && 
b[33347] == 33347 && 
b[33348] == 33348 && 
b[33349] == 33349 && 
b[33350] == 33350 && 
b[33351] == 33351 && 
b[33352] == 33352 && 
b[33353] == 33353 && 
b[33354] == 33354 && 
b[33355] == 33355 && 
b[33356] == 33356 && 
b[33357] == 33357 && 
b[33358] == 33358 && 
b[33359] == 33359 && 
b[33360] == 33360 && 
b[33361] == 33361 && 
b[33362] == 33362 && 
b[33363] == 33363 && 
b[33364] == 33364 && 
b[33365] == 33365 && 
b[33366] == 33366 && 
b[33367] == 33367 && 
b[33368] == 33368 && 
b[33369] == 33369 && 
b[33370] == 33370 && 
b[33371] == 33371 && 
b[33372] == 33372 && 
b[33373] == 33373 && 
b[33374] == 33374 && 
b[33375] == 33375 && 
b[33376] == 33376 && 
b[33377] == 33377 && 
b[33378] == 33378 && 
b[33379] == 33379 && 
b[33380] == 33380 && 
b[33381] == 33381 && 
b[33382] == 33382 && 
b[33383] == 33383 && 
b[33384] == 33384 && 
b[33385] == 33385 && 
b[33386] == 33386 && 
b[33387] == 33387 && 
b[33388] == 33388 && 
b[33389] == 33389 && 
b[33390] == 33390 && 
b[33391] == 33391 && 
b[33392] == 33392 && 
b[33393] == 33393 && 
b[33394] == 33394 && 
b[33395] == 33395 && 
b[33396] == 33396 && 
b[33397] == 33397 && 
b[33398] == 33398 && 
b[33399] == 33399 && 
b[33400] == 33400 && 
b[33401] == 33401 && 
b[33402] == 33402 && 
b[33403] == 33403 && 
b[33404] == 33404 && 
b[33405] == 33405 && 
b[33406] == 33406 && 
b[33407] == 33407 && 
b[33408] == 33408 && 
b[33409] == 33409 && 
b[33410] == 33410 && 
b[33411] == 33411 && 
b[33412] == 33412 && 
b[33413] == 33413 && 
b[33414] == 33414 && 
b[33415] == 33415 && 
b[33416] == 33416 && 
b[33417] == 33417 && 
b[33418] == 33418 && 
b[33419] == 33419 && 
b[33420] == 33420 && 
b[33421] == 33421 && 
b[33422] == 33422 && 
b[33423] == 33423 && 
b[33424] == 33424 && 
b[33425] == 33425 && 
b[33426] == 33426 && 
b[33427] == 33427 && 
b[33428] == 33428 && 
b[33429] == 33429 && 
b[33430] == 33430 && 
b[33431] == 33431 && 
b[33432] == 33432 && 
b[33433] == 33433 && 
b[33434] == 33434 && 
b[33435] == 33435 && 
b[33436] == 33436 && 
b[33437] == 33437 && 
b[33438] == 33438 && 
b[33439] == 33439 && 
b[33440] == 33440 && 
b[33441] == 33441 && 
b[33442] == 33442 && 
b[33443] == 33443 && 
b[33444] == 33444 && 
b[33445] == 33445 && 
b[33446] == 33446 && 
b[33447] == 33447 && 
b[33448] == 33448 && 
b[33449] == 33449 && 
b[33450] == 33450 && 
b[33451] == 33451 && 
b[33452] == 33452 && 
b[33453] == 33453 && 
b[33454] == 33454 && 
b[33455] == 33455 && 
b[33456] == 33456 && 
b[33457] == 33457 && 
b[33458] == 33458 && 
b[33459] == 33459 && 
b[33460] == 33460 && 
b[33461] == 33461 && 
b[33462] == 33462 && 
b[33463] == 33463 && 
b[33464] == 33464 && 
b[33465] == 33465 && 
b[33466] == 33466 && 
b[33467] == 33467 && 
b[33468] == 33468 && 
b[33469] == 33469 && 
b[33470] == 33470 && 
b[33471] == 33471 && 
b[33472] == 33472 && 
b[33473] == 33473 && 
b[33474] == 33474 && 
b[33475] == 33475 && 
b[33476] == 33476 && 
b[33477] == 33477 && 
b[33478] == 33478 && 
b[33479] == 33479 && 
b[33480] == 33480 && 
b[33481] == 33481 && 
b[33482] == 33482 && 
b[33483] == 33483 && 
b[33484] == 33484 && 
b[33485] == 33485 && 
b[33486] == 33486 && 
b[33487] == 33487 && 
b[33488] == 33488 && 
b[33489] == 33489 && 
b[33490] == 33490 && 
b[33491] == 33491 && 
b[33492] == 33492 && 
b[33493] == 33493 && 
b[33494] == 33494 && 
b[33495] == 33495 && 
b[33496] == 33496 && 
b[33497] == 33497 && 
b[33498] == 33498 && 
b[33499] == 33499 && 
b[33500] == 33500 && 
b[33501] == 33501 && 
b[33502] == 33502 && 
b[33503] == 33503 && 
b[33504] == 33504 && 
b[33505] == 33505 && 
b[33506] == 33506 && 
b[33507] == 33507 && 
b[33508] == 33508 && 
b[33509] == 33509 && 
b[33510] == 33510 && 
b[33511] == 33511 && 
b[33512] == 33512 && 
b[33513] == 33513 && 
b[33514] == 33514 && 
b[33515] == 33515 && 
b[33516] == 33516 && 
b[33517] == 33517 && 
b[33518] == 33518 && 
b[33519] == 33519 && 
b[33520] == 33520 && 
b[33521] == 33521 && 
b[33522] == 33522 && 
b[33523] == 33523 && 
b[33524] == 33524 && 
b[33525] == 33525 && 
b[33526] == 33526 && 
b[33527] == 33527 && 
b[33528] == 33528 && 
b[33529] == 33529 && 
b[33530] == 33530 && 
b[33531] == 33531 && 
b[33532] == 33532 && 
b[33533] == 33533 && 
b[33534] == 33534 && 
b[33535] == 33535 && 
b[33536] == 33536 && 
b[33537] == 33537 && 
b[33538] == 33538 && 
b[33539] == 33539 && 
b[33540] == 33540 && 
b[33541] == 33541 && 
b[33542] == 33542 && 
b[33543] == 33543 && 
b[33544] == 33544 && 
b[33545] == 33545 && 
b[33546] == 33546 && 
b[33547] == 33547 && 
b[33548] == 33548 && 
b[33549] == 33549 && 
b[33550] == 33550 && 
b[33551] == 33551 && 
b[33552] == 33552 && 
b[33553] == 33553 && 
b[33554] == 33554 && 
b[33555] == 33555 && 
b[33556] == 33556 && 
b[33557] == 33557 && 
b[33558] == 33558 && 
b[33559] == 33559 && 
b[33560] == 33560 && 
b[33561] == 33561 && 
b[33562] == 33562 && 
b[33563] == 33563 && 
b[33564] == 33564 && 
b[33565] == 33565 && 
b[33566] == 33566 && 
b[33567] == 33567 && 
b[33568] == 33568 && 
b[33569] == 33569 && 
b[33570] == 33570 && 
b[33571] == 33571 && 
b[33572] == 33572 && 
b[33573] == 33573 && 
b[33574] == 33574 && 
b[33575] == 33575 && 
b[33576] == 33576 && 
b[33577] == 33577 && 
b[33578] == 33578 && 
b[33579] == 33579 && 
b[33580] == 33580 && 
b[33581] == 33581 && 
b[33582] == 33582 && 
b[33583] == 33583 && 
b[33584] == 33584 && 
b[33585] == 33585 && 
b[33586] == 33586 && 
b[33587] == 33587 && 
b[33588] == 33588 && 
b[33589] == 33589 && 
b[33590] == 33590 && 
b[33591] == 33591 && 
b[33592] == 33592 && 
b[33593] == 33593 && 
b[33594] == 33594 && 
b[33595] == 33595 && 
b[33596] == 33596 && 
b[33597] == 33597 && 
b[33598] == 33598 && 
b[33599] == 33599 && 
b[33600] == 33600 && 
b[33601] == 33601 && 
b[33602] == 33602 && 
b[33603] == 33603 && 
b[33604] == 33604 && 
b[33605] == 33605 && 
b[33606] == 33606 && 
b[33607] == 33607 && 
b[33608] == 33608 && 
b[33609] == 33609 && 
b[33610] == 33610 && 
b[33611] == 33611 && 
b[33612] == 33612 && 
b[33613] == 33613 && 
b[33614] == 33614 && 
b[33615] == 33615 && 
b[33616] == 33616 && 
b[33617] == 33617 && 
b[33618] == 33618 && 
b[33619] == 33619 && 
b[33620] == 33620 && 
b[33621] == 33621 && 
b[33622] == 33622 && 
b[33623] == 33623 && 
b[33624] == 33624 && 
b[33625] == 33625 && 
b[33626] == 33626 && 
b[33627] == 33627 && 
b[33628] == 33628 && 
b[33629] == 33629 && 
b[33630] == 33630 && 
b[33631] == 33631 && 
b[33632] == 33632 && 
b[33633] == 33633 && 
b[33634] == 33634 && 
b[33635] == 33635 && 
b[33636] == 33636 && 
b[33637] == 33637 && 
b[33638] == 33638 && 
b[33639] == 33639 && 
b[33640] == 33640 && 
b[33641] == 33641 && 
b[33642] == 33642 && 
b[33643] == 33643 && 
b[33644] == 33644 && 
b[33645] == 33645 && 
b[33646] == 33646 && 
b[33647] == 33647 && 
b[33648] == 33648 && 
b[33649] == 33649 && 
b[33650] == 33650 && 
b[33651] == 33651 && 
b[33652] == 33652 && 
b[33653] == 33653 && 
b[33654] == 33654 && 
b[33655] == 33655 && 
b[33656] == 33656 && 
b[33657] == 33657 && 
b[33658] == 33658 && 
b[33659] == 33659 && 
b[33660] == 33660 && 
b[33661] == 33661 && 
b[33662] == 33662 && 
b[33663] == 33663 && 
b[33664] == 33664 && 
b[33665] == 33665 && 
b[33666] == 33666 && 
b[33667] == 33667 && 
b[33668] == 33668 && 
b[33669] == 33669 && 
b[33670] == 33670 && 
b[33671] == 33671 && 
b[33672] == 33672 && 
b[33673] == 33673 && 
b[33674] == 33674 && 
b[33675] == 33675 && 
b[33676] == 33676 && 
b[33677] == 33677 && 
b[33678] == 33678 && 
b[33679] == 33679 && 
b[33680] == 33680 && 
b[33681] == 33681 && 
b[33682] == 33682 && 
b[33683] == 33683 && 
b[33684] == 33684 && 
b[33685] == 33685 && 
b[33686] == 33686 && 
b[33687] == 33687 && 
b[33688] == 33688 && 
b[33689] == 33689 && 
b[33690] == 33690 && 
b[33691] == 33691 && 
b[33692] == 33692 && 
b[33693] == 33693 && 
b[33694] == 33694 && 
b[33695] == 33695 && 
b[33696] == 33696 && 
b[33697] == 33697 && 
b[33698] == 33698 && 
b[33699] == 33699 && 
b[33700] == 33700 && 
b[33701] == 33701 && 
b[33702] == 33702 && 
b[33703] == 33703 && 
b[33704] == 33704 && 
b[33705] == 33705 && 
b[33706] == 33706 && 
b[33707] == 33707 && 
b[33708] == 33708 && 
b[33709] == 33709 && 
b[33710] == 33710 && 
b[33711] == 33711 && 
b[33712] == 33712 && 
b[33713] == 33713 && 
b[33714] == 33714 && 
b[33715] == 33715 && 
b[33716] == 33716 && 
b[33717] == 33717 && 
b[33718] == 33718 && 
b[33719] == 33719 && 
b[33720] == 33720 && 
b[33721] == 33721 && 
b[33722] == 33722 && 
b[33723] == 33723 && 
b[33724] == 33724 && 
b[33725] == 33725 && 
b[33726] == 33726 && 
b[33727] == 33727 && 
b[33728] == 33728 && 
b[33729] == 33729 && 
b[33730] == 33730 && 
b[33731] == 33731 && 
b[33732] == 33732 && 
b[33733] == 33733 && 
b[33734] == 33734 && 
b[33735] == 33735 && 
b[33736] == 33736 && 
b[33737] == 33737 && 
b[33738] == 33738 && 
b[33739] == 33739 && 
b[33740] == 33740 && 
b[33741] == 33741 && 
b[33742] == 33742 && 
b[33743] == 33743 && 
b[33744] == 33744 && 
b[33745] == 33745 && 
b[33746] == 33746 && 
b[33747] == 33747 && 
b[33748] == 33748 && 
b[33749] == 33749 && 
b[33750] == 33750 && 
b[33751] == 33751 && 
b[33752] == 33752 && 
b[33753] == 33753 && 
b[33754] == 33754 && 
b[33755] == 33755 && 
b[33756] == 33756 && 
b[33757] == 33757 && 
b[33758] == 33758 && 
b[33759] == 33759 && 
b[33760] == 33760 && 
b[33761] == 33761 && 
b[33762] == 33762 && 
b[33763] == 33763 && 
b[33764] == 33764 && 
b[33765] == 33765 && 
b[33766] == 33766 && 
b[33767] == 33767 && 
b[33768] == 33768 && 
b[33769] == 33769 && 
b[33770] == 33770 && 
b[33771] == 33771 && 
b[33772] == 33772 && 
b[33773] == 33773 && 
b[33774] == 33774 && 
b[33775] == 33775 && 
b[33776] == 33776 && 
b[33777] == 33777 && 
b[33778] == 33778 && 
b[33779] == 33779 && 
b[33780] == 33780 && 
b[33781] == 33781 && 
b[33782] == 33782 && 
b[33783] == 33783 && 
b[33784] == 33784 && 
b[33785] == 33785 && 
b[33786] == 33786 && 
b[33787] == 33787 && 
b[33788] == 33788 && 
b[33789] == 33789 && 
b[33790] == 33790 && 
b[33791] == 33791 && 
b[33792] == 33792 && 
b[33793] == 33793 && 
b[33794] == 33794 && 
b[33795] == 33795 && 
b[33796] == 33796 && 
b[33797] == 33797 && 
b[33798] == 33798 && 
b[33799] == 33799 && 
b[33800] == 33800 && 
b[33801] == 33801 && 
b[33802] == 33802 && 
b[33803] == 33803 && 
b[33804] == 33804 && 
b[33805] == 33805 && 
b[33806] == 33806 && 
b[33807] == 33807 && 
b[33808] == 33808 && 
b[33809] == 33809 && 
b[33810] == 33810 && 
b[33811] == 33811 && 
b[33812] == 33812 && 
b[33813] == 33813 && 
b[33814] == 33814 && 
b[33815] == 33815 && 
b[33816] == 33816 && 
b[33817] == 33817 && 
b[33818] == 33818 && 
b[33819] == 33819 && 
b[33820] == 33820 && 
b[33821] == 33821 && 
b[33822] == 33822 && 
b[33823] == 33823 && 
b[33824] == 33824 && 
b[33825] == 33825 && 
b[33826] == 33826 && 
b[33827] == 33827 && 
b[33828] == 33828 && 
b[33829] == 33829 && 
b[33830] == 33830 && 
b[33831] == 33831 && 
b[33832] == 33832 && 
b[33833] == 33833 && 
b[33834] == 33834 && 
b[33835] == 33835 && 
b[33836] == 33836 && 
b[33837] == 33837 && 
b[33838] == 33838 && 
b[33839] == 33839 && 
b[33840] == 33840 && 
b[33841] == 33841 && 
b[33842] == 33842 && 
b[33843] == 33843 && 
b[33844] == 33844 && 
b[33845] == 33845 && 
b[33846] == 33846 && 
b[33847] == 33847 && 
b[33848] == 33848 && 
b[33849] == 33849 && 
b[33850] == 33850 && 
b[33851] == 33851 && 
b[33852] == 33852 && 
b[33853] == 33853 && 
b[33854] == 33854 && 
b[33855] == 33855 && 
b[33856] == 33856 && 
b[33857] == 33857 && 
b[33858] == 33858 && 
b[33859] == 33859 && 
b[33860] == 33860 && 
b[33861] == 33861 && 
b[33862] == 33862 && 
b[33863] == 33863 && 
b[33864] == 33864 && 
b[33865] == 33865 && 
b[33866] == 33866 && 
b[33867] == 33867 && 
b[33868] == 33868 && 
b[33869] == 33869 && 
b[33870] == 33870 && 
b[33871] == 33871 && 
b[33872] == 33872 && 
b[33873] == 33873 && 
b[33874] == 33874 && 
b[33875] == 33875 && 
b[33876] == 33876 && 
b[33877] == 33877 && 
b[33878] == 33878 && 
b[33879] == 33879 && 
b[33880] == 33880 && 
b[33881] == 33881 && 
b[33882] == 33882 && 
b[33883] == 33883 && 
b[33884] == 33884 && 
b[33885] == 33885 && 
b[33886] == 33886 && 
b[33887] == 33887 && 
b[33888] == 33888 && 
b[33889] == 33889 && 
b[33890] == 33890 && 
b[33891] == 33891 && 
b[33892] == 33892 && 
b[33893] == 33893 && 
b[33894] == 33894 && 
b[33895] == 33895 && 
b[33896] == 33896 && 
b[33897] == 33897 && 
b[33898] == 33898 && 
b[33899] == 33899 && 
b[33900] == 33900 && 
b[33901] == 33901 && 
b[33902] == 33902 && 
b[33903] == 33903 && 
b[33904] == 33904 && 
b[33905] == 33905 && 
b[33906] == 33906 && 
b[33907] == 33907 && 
b[33908] == 33908 && 
b[33909] == 33909 && 
b[33910] == 33910 && 
b[33911] == 33911 && 
b[33912] == 33912 && 
b[33913] == 33913 && 
b[33914] == 33914 && 
b[33915] == 33915 && 
b[33916] == 33916 && 
b[33917] == 33917 && 
b[33918] == 33918 && 
b[33919] == 33919 && 
b[33920] == 33920 && 
b[33921] == 33921 && 
b[33922] == 33922 && 
b[33923] == 33923 && 
b[33924] == 33924 && 
b[33925] == 33925 && 
b[33926] == 33926 && 
b[33927] == 33927 && 
b[33928] == 33928 && 
b[33929] == 33929 && 
b[33930] == 33930 && 
b[33931] == 33931 && 
b[33932] == 33932 && 
b[33933] == 33933 && 
b[33934] == 33934 && 
b[33935] == 33935 && 
b[33936] == 33936 && 
b[33937] == 33937 && 
b[33938] == 33938 && 
b[33939] == 33939 && 
b[33940] == 33940 && 
b[33941] == 33941 && 
b[33942] == 33942 && 
b[33943] == 33943 && 
b[33944] == 33944 && 
b[33945] == 33945 && 
b[33946] == 33946 && 
b[33947] == 33947 && 
b[33948] == 33948 && 
b[33949] == 33949 && 
b[33950] == 33950 && 
b[33951] == 33951 && 
b[33952] == 33952 && 
b[33953] == 33953 && 
b[33954] == 33954 && 
b[33955] == 33955 && 
b[33956] == 33956 && 
b[33957] == 33957 && 
b[33958] == 33958 && 
b[33959] == 33959 && 
b[33960] == 33960 && 
b[33961] == 33961 && 
b[33962] == 33962 && 
b[33963] == 33963 && 
b[33964] == 33964 && 
b[33965] == 33965 && 
b[33966] == 33966 && 
b[33967] == 33967 && 
b[33968] == 33968 && 
b[33969] == 33969 && 
b[33970] == 33970 && 
b[33971] == 33971 && 
b[33972] == 33972 && 
b[33973] == 33973 && 
b[33974] == 33974 && 
b[33975] == 33975 && 
b[33976] == 33976 && 
b[33977] == 33977 && 
b[33978] == 33978 && 
b[33979] == 33979 && 
b[33980] == 33980 && 
b[33981] == 33981 && 
b[33982] == 33982 && 
b[33983] == 33983 && 
b[33984] == 33984 && 
b[33985] == 33985 && 
b[33986] == 33986 && 
b[33987] == 33987 && 
b[33988] == 33988 && 
b[33989] == 33989 && 
b[33990] == 33990 && 
b[33991] == 33991 && 
b[33992] == 33992 && 
b[33993] == 33993 && 
b[33994] == 33994 && 
b[33995] == 33995 && 
b[33996] == 33996 && 
b[33997] == 33997 && 
b[33998] == 33998 && 
b[33999] == 33999 && 
b[34000] == 34000 && 
b[34001] == 34001 && 
b[34002] == 34002 && 
b[34003] == 34003 && 
b[34004] == 34004 && 
b[34005] == 34005 && 
b[34006] == 34006 && 
b[34007] == 34007 && 
b[34008] == 34008 && 
b[34009] == 34009 && 
b[34010] == 34010 && 
b[34011] == 34011 && 
b[34012] == 34012 && 
b[34013] == 34013 && 
b[34014] == 34014 && 
b[34015] == 34015 && 
b[34016] == 34016 && 
b[34017] == 34017 && 
b[34018] == 34018 && 
b[34019] == 34019 && 
b[34020] == 34020 && 
b[34021] == 34021 && 
b[34022] == 34022 && 
b[34023] == 34023 && 
b[34024] == 34024 && 
b[34025] == 34025 && 
b[34026] == 34026 && 
b[34027] == 34027 && 
b[34028] == 34028 && 
b[34029] == 34029 && 
b[34030] == 34030 && 
b[34031] == 34031 && 
b[34032] == 34032 && 
b[34033] == 34033 && 
b[34034] == 34034 && 
b[34035] == 34035 && 
b[34036] == 34036 && 
b[34037] == 34037 && 
b[34038] == 34038 && 
b[34039] == 34039 && 
b[34040] == 34040 && 
b[34041] == 34041 && 
b[34042] == 34042 && 
b[34043] == 34043 && 
b[34044] == 34044 && 
b[34045] == 34045 && 
b[34046] == 34046 && 
b[34047] == 34047 && 
b[34048] == 34048 && 
b[34049] == 34049 && 
b[34050] == 34050 && 
b[34051] == 34051 && 
b[34052] == 34052 && 
b[34053] == 34053 && 
b[34054] == 34054 && 
b[34055] == 34055 && 
b[34056] == 34056 && 
b[34057] == 34057 && 
b[34058] == 34058 && 
b[34059] == 34059 && 
b[34060] == 34060 && 
b[34061] == 34061 && 
b[34062] == 34062 && 
b[34063] == 34063 && 
b[34064] == 34064 && 
b[34065] == 34065 && 
b[34066] == 34066 && 
b[34067] == 34067 && 
b[34068] == 34068 && 
b[34069] == 34069 && 
b[34070] == 34070 && 
b[34071] == 34071 && 
b[34072] == 34072 && 
b[34073] == 34073 && 
b[34074] == 34074 && 
b[34075] == 34075 && 
b[34076] == 34076 && 
b[34077] == 34077 && 
b[34078] == 34078 && 
b[34079] == 34079 && 
b[34080] == 34080 && 
b[34081] == 34081 && 
b[34082] == 34082 && 
b[34083] == 34083 && 
b[34084] == 34084 && 
b[34085] == 34085 && 
b[34086] == 34086 && 
b[34087] == 34087 && 
b[34088] == 34088 && 
b[34089] == 34089 && 
b[34090] == 34090 && 
b[34091] == 34091 && 
b[34092] == 34092 && 
b[34093] == 34093 && 
b[34094] == 34094 && 
b[34095] == 34095 && 
b[34096] == 34096 && 
b[34097] == 34097 && 
b[34098] == 34098 && 
b[34099] == 34099 && 
b[34100] == 34100 && 
b[34101] == 34101 && 
b[34102] == 34102 && 
b[34103] == 34103 && 
b[34104] == 34104 && 
b[34105] == 34105 && 
b[34106] == 34106 && 
b[34107] == 34107 && 
b[34108] == 34108 && 
b[34109] == 34109 && 
b[34110] == 34110 && 
b[34111] == 34111 && 
b[34112] == 34112 && 
b[34113] == 34113 && 
b[34114] == 34114 && 
b[34115] == 34115 && 
b[34116] == 34116 && 
b[34117] == 34117 && 
b[34118] == 34118 && 
b[34119] == 34119 && 
b[34120] == 34120 && 
b[34121] == 34121 && 
b[34122] == 34122 && 
b[34123] == 34123 && 
b[34124] == 34124 && 
b[34125] == 34125 && 
b[34126] == 34126 && 
b[34127] == 34127 && 
b[34128] == 34128 && 
b[34129] == 34129 && 
b[34130] == 34130 && 
b[34131] == 34131 && 
b[34132] == 34132 && 
b[34133] == 34133 && 
b[34134] == 34134 && 
b[34135] == 34135 && 
b[34136] == 34136 && 
b[34137] == 34137 && 
b[34138] == 34138 && 
b[34139] == 34139 && 
b[34140] == 34140 && 
b[34141] == 34141 && 
b[34142] == 34142 && 
b[34143] == 34143 && 
b[34144] == 34144 && 
b[34145] == 34145 && 
b[34146] == 34146 && 
b[34147] == 34147 && 
b[34148] == 34148 && 
b[34149] == 34149 && 
b[34150] == 34150 && 
b[34151] == 34151 && 
b[34152] == 34152 && 
b[34153] == 34153 && 
b[34154] == 34154 && 
b[34155] == 34155 && 
b[34156] == 34156 && 
b[34157] == 34157 && 
b[34158] == 34158 && 
b[34159] == 34159 && 
b[34160] == 34160 && 
b[34161] == 34161 && 
b[34162] == 34162 && 
b[34163] == 34163 && 
b[34164] == 34164 && 
b[34165] == 34165 && 
b[34166] == 34166 && 
b[34167] == 34167 && 
b[34168] == 34168 && 
b[34169] == 34169 && 
b[34170] == 34170 && 
b[34171] == 34171 && 
b[34172] == 34172 && 
b[34173] == 34173 && 
b[34174] == 34174 && 
b[34175] == 34175 && 
b[34176] == 34176 && 
b[34177] == 34177 && 
b[34178] == 34178 && 
b[34179] == 34179 && 
b[34180] == 34180 && 
b[34181] == 34181 && 
b[34182] == 34182 && 
b[34183] == 34183 && 
b[34184] == 34184 && 
b[34185] == 34185 && 
b[34186] == 34186 && 
b[34187] == 34187 && 
b[34188] == 34188 && 
b[34189] == 34189 && 
b[34190] == 34190 && 
b[34191] == 34191 && 
b[34192] == 34192 && 
b[34193] == 34193 && 
b[34194] == 34194 && 
b[34195] == 34195 && 
b[34196] == 34196 && 
b[34197] == 34197 && 
b[34198] == 34198 && 
b[34199] == 34199 && 
b[34200] == 34200 && 
b[34201] == 34201 && 
b[34202] == 34202 && 
b[34203] == 34203 && 
b[34204] == 34204 && 
b[34205] == 34205 && 
b[34206] == 34206 && 
b[34207] == 34207 && 
b[34208] == 34208 && 
b[34209] == 34209 && 
b[34210] == 34210 && 
b[34211] == 34211 && 
b[34212] == 34212 && 
b[34213] == 34213 && 
b[34214] == 34214 && 
b[34215] == 34215 && 
b[34216] == 34216 && 
b[34217] == 34217 && 
b[34218] == 34218 && 
b[34219] == 34219 && 
b[34220] == 34220 && 
b[34221] == 34221 && 
b[34222] == 34222 && 
b[34223] == 34223 && 
b[34224] == 34224 && 
b[34225] == 34225 && 
b[34226] == 34226 && 
b[34227] == 34227 && 
b[34228] == 34228 && 
b[34229] == 34229 && 
b[34230] == 34230 && 
b[34231] == 34231 && 
b[34232] == 34232 && 
b[34233] == 34233 && 
b[34234] == 34234 && 
b[34235] == 34235 && 
b[34236] == 34236 && 
b[34237] == 34237 && 
b[34238] == 34238 && 
b[34239] == 34239 && 
b[34240] == 34240 && 
b[34241] == 34241 && 
b[34242] == 34242 && 
b[34243] == 34243 && 
b[34244] == 34244 && 
b[34245] == 34245 && 
b[34246] == 34246 && 
b[34247] == 34247 && 
b[34248] == 34248 && 
b[34249] == 34249 && 
b[34250] == 34250 && 
b[34251] == 34251 && 
b[34252] == 34252 && 
b[34253] == 34253 && 
b[34254] == 34254 && 
b[34255] == 34255 && 
b[34256] == 34256 && 
b[34257] == 34257 && 
b[34258] == 34258 && 
b[34259] == 34259 && 
b[34260] == 34260 && 
b[34261] == 34261 && 
b[34262] == 34262 && 
b[34263] == 34263 && 
b[34264] == 34264 && 
b[34265] == 34265 && 
b[34266] == 34266 && 
b[34267] == 34267 && 
b[34268] == 34268 && 
b[34269] == 34269 && 
b[34270] == 34270 && 
b[34271] == 34271 && 
b[34272] == 34272 && 
b[34273] == 34273 && 
b[34274] == 34274 && 
b[34275] == 34275 && 
b[34276] == 34276 && 
b[34277] == 34277 && 
b[34278] == 34278 && 
b[34279] == 34279 && 
b[34280] == 34280 && 
b[34281] == 34281 && 
b[34282] == 34282 && 
b[34283] == 34283 && 
b[34284] == 34284 && 
b[34285] == 34285 && 
b[34286] == 34286 && 
b[34287] == 34287 && 
b[34288] == 34288 && 
b[34289] == 34289 && 
b[34290] == 34290 && 
b[34291] == 34291 && 
b[34292] == 34292 && 
b[34293] == 34293 && 
b[34294] == 34294 && 
b[34295] == 34295 && 
b[34296] == 34296 && 
b[34297] == 34297 && 
b[34298] == 34298 && 
b[34299] == 34299 && 
b[34300] == 34300 && 
b[34301] == 34301 && 
b[34302] == 34302 && 
b[34303] == 34303 && 
b[34304] == 34304 && 
b[34305] == 34305 && 
b[34306] == 34306 && 
b[34307] == 34307 && 
b[34308] == 34308 && 
b[34309] == 34309 && 
b[34310] == 34310 && 
b[34311] == 34311 && 
b[34312] == 34312 && 
b[34313] == 34313 && 
b[34314] == 34314 && 
b[34315] == 34315 && 
b[34316] == 34316 && 
b[34317] == 34317 && 
b[34318] == 34318 && 
b[34319] == 34319 && 
b[34320] == 34320 && 
b[34321] == 34321 && 
b[34322] == 34322 && 
b[34323] == 34323 && 
b[34324] == 34324 && 
b[34325] == 34325 && 
b[34326] == 34326 && 
b[34327] == 34327 && 
b[34328] == 34328 && 
b[34329] == 34329 && 
b[34330] == 34330 && 
b[34331] == 34331 && 
b[34332] == 34332 && 
b[34333] == 34333 && 
b[34334] == 34334 && 
b[34335] == 34335 && 
b[34336] == 34336 && 
b[34337] == 34337 && 
b[34338] == 34338 && 
b[34339] == 34339 && 
b[34340] == 34340 && 
b[34341] == 34341 && 
b[34342] == 34342 && 
b[34343] == 34343 && 
b[34344] == 34344 && 
b[34345] == 34345 && 
b[34346] == 34346 && 
b[34347] == 34347 && 
b[34348] == 34348 && 
b[34349] == 34349 && 
b[34350] == 34350 && 
b[34351] == 34351 && 
b[34352] == 34352 && 
b[34353] == 34353 && 
b[34354] == 34354 && 
b[34355] == 34355 && 
b[34356] == 34356 && 
b[34357] == 34357 && 
b[34358] == 34358 && 
b[34359] == 34359 && 
b[34360] == 34360 && 
b[34361] == 34361 && 
b[34362] == 34362 && 
b[34363] == 34363 && 
b[34364] == 34364 && 
b[34365] == 34365 && 
b[34366] == 34366 && 
b[34367] == 34367 && 
b[34368] == 34368 && 
b[34369] == 34369 && 
b[34370] == 34370 && 
b[34371] == 34371 && 
b[34372] == 34372 && 
b[34373] == 34373 && 
b[34374] == 34374 && 
b[34375] == 34375 && 
b[34376] == 34376 && 
b[34377] == 34377 && 
b[34378] == 34378 && 
b[34379] == 34379 && 
b[34380] == 34380 && 
b[34381] == 34381 && 
b[34382] == 34382 && 
b[34383] == 34383 && 
b[34384] == 34384 && 
b[34385] == 34385 && 
b[34386] == 34386 && 
b[34387] == 34387 && 
b[34388] == 34388 && 
b[34389] == 34389 && 
b[34390] == 34390 && 
b[34391] == 34391 && 
b[34392] == 34392 && 
b[34393] == 34393 && 
b[34394] == 34394 && 
b[34395] == 34395 && 
b[34396] == 34396 && 
b[34397] == 34397 && 
b[34398] == 34398 && 
b[34399] == 34399 && 
b[34400] == 34400 && 
b[34401] == 34401 && 
b[34402] == 34402 && 
b[34403] == 34403 && 
b[34404] == 34404 && 
b[34405] == 34405 && 
b[34406] == 34406 && 
b[34407] == 34407 && 
b[34408] == 34408 && 
b[34409] == 34409 && 
b[34410] == 34410 && 
b[34411] == 34411 && 
b[34412] == 34412 && 
b[34413] == 34413 && 
b[34414] == 34414 && 
b[34415] == 34415 && 
b[34416] == 34416 && 
b[34417] == 34417 && 
b[34418] == 34418 && 
b[34419] == 34419 && 
b[34420] == 34420 && 
b[34421] == 34421 && 
b[34422] == 34422 && 
b[34423] == 34423 && 
b[34424] == 34424 && 
b[34425] == 34425 && 
b[34426] == 34426 && 
b[34427] == 34427 && 
b[34428] == 34428 && 
b[34429] == 34429 && 
b[34430] == 34430 && 
b[34431] == 34431 && 
b[34432] == 34432 && 
b[34433] == 34433 && 
b[34434] == 34434 && 
b[34435] == 34435 && 
b[34436] == 34436 && 
b[34437] == 34437 && 
b[34438] == 34438 && 
b[34439] == 34439 && 
b[34440] == 34440 && 
b[34441] == 34441 && 
b[34442] == 34442 && 
b[34443] == 34443 && 
b[34444] == 34444 && 
b[34445] == 34445 && 
b[34446] == 34446 && 
b[34447] == 34447 && 
b[34448] == 34448 && 
b[34449] == 34449 && 
b[34450] == 34450 && 
b[34451] == 34451 && 
b[34452] == 34452 && 
b[34453] == 34453 && 
b[34454] == 34454 && 
b[34455] == 34455 && 
b[34456] == 34456 && 
b[34457] == 34457 && 
b[34458] == 34458 && 
b[34459] == 34459 && 
b[34460] == 34460 && 
b[34461] == 34461 && 
b[34462] == 34462 && 
b[34463] == 34463 && 
b[34464] == 34464 && 
b[34465] == 34465 && 
b[34466] == 34466 && 
b[34467] == 34467 && 
b[34468] == 34468 && 
b[34469] == 34469 && 
b[34470] == 34470 && 
b[34471] == 34471 && 
b[34472] == 34472 && 
b[34473] == 34473 && 
b[34474] == 34474 && 
b[34475] == 34475 && 
b[34476] == 34476 && 
b[34477] == 34477 && 
b[34478] == 34478 && 
b[34479] == 34479 && 
b[34480] == 34480 && 
b[34481] == 34481 && 
b[34482] == 34482 && 
b[34483] == 34483 && 
b[34484] == 34484 && 
b[34485] == 34485 && 
b[34486] == 34486 && 
b[34487] == 34487 && 
b[34488] == 34488 && 
b[34489] == 34489 && 
b[34490] == 34490 && 
b[34491] == 34491 && 
b[34492] == 34492 && 
b[34493] == 34493 && 
b[34494] == 34494 && 
b[34495] == 34495 && 
b[34496] == 34496 && 
b[34497] == 34497 && 
b[34498] == 34498 && 
b[34499] == 34499 && 
b[34500] == 34500 && 
b[34501] == 34501 && 
b[34502] == 34502 && 
b[34503] == 34503 && 
b[34504] == 34504 && 
b[34505] == 34505 && 
b[34506] == 34506 && 
b[34507] == 34507 && 
b[34508] == 34508 && 
b[34509] == 34509 && 
b[34510] == 34510 && 
b[34511] == 34511 && 
b[34512] == 34512 && 
b[34513] == 34513 && 
b[34514] == 34514 && 
b[34515] == 34515 && 
b[34516] == 34516 && 
b[34517] == 34517 && 
b[34518] == 34518 && 
b[34519] == 34519 && 
b[34520] == 34520 && 
b[34521] == 34521 && 
b[34522] == 34522 && 
b[34523] == 34523 && 
b[34524] == 34524 && 
b[34525] == 34525 && 
b[34526] == 34526 && 
b[34527] == 34527 && 
b[34528] == 34528 && 
b[34529] == 34529 && 
b[34530] == 34530 && 
b[34531] == 34531 && 
b[34532] == 34532 && 
b[34533] == 34533 && 
b[34534] == 34534 && 
b[34535] == 34535 && 
b[34536] == 34536 && 
b[34537] == 34537 && 
b[34538] == 34538 && 
b[34539] == 34539 && 
b[34540] == 34540 && 
b[34541] == 34541 && 
b[34542] == 34542 && 
b[34543] == 34543 && 
b[34544] == 34544 && 
b[34545] == 34545 && 
b[34546] == 34546 && 
b[34547] == 34547 && 
b[34548] == 34548 && 
b[34549] == 34549 && 
b[34550] == 34550 && 
b[34551] == 34551 && 
b[34552] == 34552 && 
b[34553] == 34553 && 
b[34554] == 34554 && 
b[34555] == 34555 && 
b[34556] == 34556 && 
b[34557] == 34557 && 
b[34558] == 34558 && 
b[34559] == 34559 && 
b[34560] == 34560 && 
b[34561] == 34561 && 
b[34562] == 34562 && 
b[34563] == 34563 && 
b[34564] == 34564 && 
b[34565] == 34565 && 
b[34566] == 34566 && 
b[34567] == 34567 && 
b[34568] == 34568 && 
b[34569] == 34569 && 
b[34570] == 34570 && 
b[34571] == 34571 && 
b[34572] == 34572 && 
b[34573] == 34573 && 
b[34574] == 34574 && 
b[34575] == 34575 && 
b[34576] == 34576 && 
b[34577] == 34577 && 
b[34578] == 34578 && 
b[34579] == 34579 && 
b[34580] == 34580 && 
b[34581] == 34581 && 
b[34582] == 34582 && 
b[34583] == 34583 && 
b[34584] == 34584 && 
b[34585] == 34585 && 
b[34586] == 34586 && 
b[34587] == 34587 && 
b[34588] == 34588 && 
b[34589] == 34589 && 
b[34590] == 34590 && 
b[34591] == 34591 && 
b[34592] == 34592 && 
b[34593] == 34593 && 
b[34594] == 34594 && 
b[34595] == 34595 && 
b[34596] == 34596 && 
b[34597] == 34597 && 
b[34598] == 34598 && 
b[34599] == 34599 && 
b[34600] == 34600 && 
b[34601] == 34601 && 
b[34602] == 34602 && 
b[34603] == 34603 && 
b[34604] == 34604 && 
b[34605] == 34605 && 
b[34606] == 34606 && 
b[34607] == 34607 && 
b[34608] == 34608 && 
b[34609] == 34609 && 
b[34610] == 34610 && 
b[34611] == 34611 && 
b[34612] == 34612 && 
b[34613] == 34613 && 
b[34614] == 34614 && 
b[34615] == 34615 && 
b[34616] == 34616 && 
b[34617] == 34617 && 
b[34618] == 34618 && 
b[34619] == 34619 && 
b[34620] == 34620 && 
b[34621] == 34621 && 
b[34622] == 34622 && 
b[34623] == 34623 && 
b[34624] == 34624 && 
b[34625] == 34625 && 
b[34626] == 34626 && 
b[34627] == 34627 && 
b[34628] == 34628 && 
b[34629] == 34629 && 
b[34630] == 34630 && 
b[34631] == 34631 && 
b[34632] == 34632 && 
b[34633] == 34633 && 
b[34634] == 34634 && 
b[34635] == 34635 && 
b[34636] == 34636 && 
b[34637] == 34637 && 
b[34638] == 34638 && 
b[34639] == 34639 && 
b[34640] == 34640 && 
b[34641] == 34641 && 
b[34642] == 34642 && 
b[34643] == 34643 && 
b[34644] == 34644 && 
b[34645] == 34645 && 
b[34646] == 34646 && 
b[34647] == 34647 && 
b[34648] == 34648 && 
b[34649] == 34649 && 
b[34650] == 34650 && 
b[34651] == 34651 && 
b[34652] == 34652 && 
b[34653] == 34653 && 
b[34654] == 34654 && 
b[34655] == 34655 && 
b[34656] == 34656 && 
b[34657] == 34657 && 
b[34658] == 34658 && 
b[34659] == 34659 && 
b[34660] == 34660 && 
b[34661] == 34661 && 
b[34662] == 34662 && 
b[34663] == 34663 && 
b[34664] == 34664 && 
b[34665] == 34665 && 
b[34666] == 34666 && 
b[34667] == 34667 && 
b[34668] == 34668 && 
b[34669] == 34669 && 
b[34670] == 34670 && 
b[34671] == 34671 && 
b[34672] == 34672 && 
b[34673] == 34673 && 
b[34674] == 34674 && 
b[34675] == 34675 && 
b[34676] == 34676 && 
b[34677] == 34677 && 
b[34678] == 34678 && 
b[34679] == 34679 && 
b[34680] == 34680 && 
b[34681] == 34681 && 
b[34682] == 34682 && 
b[34683] == 34683 && 
b[34684] == 34684 && 
b[34685] == 34685 && 
b[34686] == 34686 && 
b[34687] == 34687 && 
b[34688] == 34688 && 
b[34689] == 34689 && 
b[34690] == 34690 && 
b[34691] == 34691 && 
b[34692] == 34692 && 
b[34693] == 34693 && 
b[34694] == 34694 && 
b[34695] == 34695 && 
b[34696] == 34696 && 
b[34697] == 34697 && 
b[34698] == 34698 && 
b[34699] == 34699 && 
b[34700] == 34700 && 
b[34701] == 34701 && 
b[34702] == 34702 && 
b[34703] == 34703 && 
b[34704] == 34704 && 
b[34705] == 34705 && 
b[34706] == 34706 && 
b[34707] == 34707 && 
b[34708] == 34708 && 
b[34709] == 34709 && 
b[34710] == 34710 && 
b[34711] == 34711 && 
b[34712] == 34712 && 
b[34713] == 34713 && 
b[34714] == 34714 && 
b[34715] == 34715 && 
b[34716] == 34716 && 
b[34717] == 34717 && 
b[34718] == 34718 && 
b[34719] == 34719 && 
b[34720] == 34720 && 
b[34721] == 34721 && 
b[34722] == 34722 && 
b[34723] == 34723 && 
b[34724] == 34724 && 
b[34725] == 34725 && 
b[34726] == 34726 && 
b[34727] == 34727 && 
b[34728] == 34728 && 
b[34729] == 34729 && 
b[34730] == 34730 && 
b[34731] == 34731 && 
b[34732] == 34732 && 
b[34733] == 34733 && 
b[34734] == 34734 && 
b[34735] == 34735 && 
b[34736] == 34736 && 
b[34737] == 34737 && 
b[34738] == 34738 && 
b[34739] == 34739 && 
b[34740] == 34740 && 
b[34741] == 34741 && 
b[34742] == 34742 && 
b[34743] == 34743 && 
b[34744] == 34744 && 
b[34745] == 34745 && 
b[34746] == 34746 && 
b[34747] == 34747 && 
b[34748] == 34748 && 
b[34749] == 34749 && 
b[34750] == 34750 && 
b[34751] == 34751 && 
b[34752] == 34752 && 
b[34753] == 34753 && 
b[34754] == 34754 && 
b[34755] == 34755 && 
b[34756] == 34756 && 
b[34757] == 34757 && 
b[34758] == 34758 && 
b[34759] == 34759 && 
b[34760] == 34760 && 
b[34761] == 34761 && 
b[34762] == 34762 && 
b[34763] == 34763 && 
b[34764] == 34764 && 
b[34765] == 34765 && 
b[34766] == 34766 && 
b[34767] == 34767 && 
b[34768] == 34768 && 
b[34769] == 34769 && 
b[34770] == 34770 && 
b[34771] == 34771 && 
b[34772] == 34772 && 
b[34773] == 34773 && 
b[34774] == 34774 && 
b[34775] == 34775 && 
b[34776] == 34776 && 
b[34777] == 34777 && 
b[34778] == 34778 && 
b[34779] == 34779 && 
b[34780] == 34780 && 
b[34781] == 34781 && 
b[34782] == 34782 && 
b[34783] == 34783 && 
b[34784] == 34784 && 
b[34785] == 34785 && 
b[34786] == 34786 && 
b[34787] == 34787 && 
b[34788] == 34788 && 
b[34789] == 34789 && 
b[34790] == 34790 && 
b[34791] == 34791 && 
b[34792] == 34792 && 
b[34793] == 34793 && 
b[34794] == 34794 && 
b[34795] == 34795 && 
b[34796] == 34796 && 
b[34797] == 34797 && 
b[34798] == 34798 && 
b[34799] == 34799 && 
b[34800] == 34800 && 
b[34801] == 34801 && 
b[34802] == 34802 && 
b[34803] == 34803 && 
b[34804] == 34804 && 
b[34805] == 34805 && 
b[34806] == 34806 && 
b[34807] == 34807 && 
b[34808] == 34808 && 
b[34809] == 34809 && 
b[34810] == 34810 && 
b[34811] == 34811 && 
b[34812] == 34812 && 
b[34813] == 34813 && 
b[34814] == 34814 && 
b[34815] == 34815 && 
b[34816] == 34816 && 
b[34817] == 34817 && 
b[34818] == 34818 && 
b[34819] == 34819 && 
b[34820] == 34820 && 
b[34821] == 34821 && 
b[34822] == 34822 && 
b[34823] == 34823 && 
b[34824] == 34824 && 
b[34825] == 34825 && 
b[34826] == 34826 && 
b[34827] == 34827 && 
b[34828] == 34828 && 
b[34829] == 34829 && 
b[34830] == 34830 && 
b[34831] == 34831 && 
b[34832] == 34832 && 
b[34833] == 34833 && 
b[34834] == 34834 && 
b[34835] == 34835 && 
b[34836] == 34836 && 
b[34837] == 34837 && 
b[34838] == 34838 && 
b[34839] == 34839 && 
b[34840] == 34840 && 
b[34841] == 34841 && 
b[34842] == 34842 && 
b[34843] == 34843 && 
b[34844] == 34844 && 
b[34845] == 34845 && 
b[34846] == 34846 && 
b[34847] == 34847 && 
b[34848] == 34848 && 
b[34849] == 34849 && 
b[34850] == 34850 && 
b[34851] == 34851 && 
b[34852] == 34852 && 
b[34853] == 34853 && 
b[34854] == 34854 && 
b[34855] == 34855 && 
b[34856] == 34856 && 
b[34857] == 34857 && 
b[34858] == 34858 && 
b[34859] == 34859 && 
b[34860] == 34860 && 
b[34861] == 34861 && 
b[34862] == 34862 && 
b[34863] == 34863 && 
b[34864] == 34864 && 
b[34865] == 34865 && 
b[34866] == 34866 && 
b[34867] == 34867 && 
b[34868] == 34868 && 
b[34869] == 34869 && 
b[34870] == 34870 && 
b[34871] == 34871 && 
b[34872] == 34872 && 
b[34873] == 34873 && 
b[34874] == 34874 && 
b[34875] == 34875 && 
b[34876] == 34876 && 
b[34877] == 34877 && 
b[34878] == 34878 && 
b[34879] == 34879 && 
b[34880] == 34880 && 
b[34881] == 34881 && 
b[34882] == 34882 && 
b[34883] == 34883 && 
b[34884] == 34884 && 
b[34885] == 34885 && 
b[34886] == 34886 && 
b[34887] == 34887 && 
b[34888] == 34888 && 
b[34889] == 34889 && 
b[34890] == 34890 && 
b[34891] == 34891 && 
b[34892] == 34892 && 
b[34893] == 34893 && 
b[34894] == 34894 && 
b[34895] == 34895 && 
b[34896] == 34896 && 
b[34897] == 34897 && 
b[34898] == 34898 && 
b[34899] == 34899 && 
b[34900] == 34900 && 
b[34901] == 34901 && 
b[34902] == 34902 && 
b[34903] == 34903 && 
b[34904] == 34904 && 
b[34905] == 34905 && 
b[34906] == 34906 && 
b[34907] == 34907 && 
b[34908] == 34908 && 
b[34909] == 34909 && 
b[34910] == 34910 && 
b[34911] == 34911 && 
b[34912] == 34912 && 
b[34913] == 34913 && 
b[34914] == 34914 && 
b[34915] == 34915 && 
b[34916] == 34916 && 
b[34917] == 34917 && 
b[34918] == 34918 && 
b[34919] == 34919 && 
b[34920] == 34920 && 
b[34921] == 34921 && 
b[34922] == 34922 && 
b[34923] == 34923 && 
b[34924] == 34924 && 
b[34925] == 34925 && 
b[34926] == 34926 && 
b[34927] == 34927 && 
b[34928] == 34928 && 
b[34929] == 34929 && 
b[34930] == 34930 && 
b[34931] == 34931 && 
b[34932] == 34932 && 
b[34933] == 34933 && 
b[34934] == 34934 && 
b[34935] == 34935 && 
b[34936] == 34936 && 
b[34937] == 34937 && 
b[34938] == 34938 && 
b[34939] == 34939 && 
b[34940] == 34940 && 
b[34941] == 34941 && 
b[34942] == 34942 && 
b[34943] == 34943 && 
b[34944] == 34944 && 
b[34945] == 34945 && 
b[34946] == 34946 && 
b[34947] == 34947 && 
b[34948] == 34948 && 
b[34949] == 34949 && 
b[34950] == 34950 && 
b[34951] == 34951 && 
b[34952] == 34952 && 
b[34953] == 34953 && 
b[34954] == 34954 && 
b[34955] == 34955 && 
b[34956] == 34956 && 
b[34957] == 34957 && 
b[34958] == 34958 && 
b[34959] == 34959 && 
b[34960] == 34960 && 
b[34961] == 34961 && 
b[34962] == 34962 && 
b[34963] == 34963 && 
b[34964] == 34964 && 
b[34965] == 34965 && 
b[34966] == 34966 && 
b[34967] == 34967 && 
b[34968] == 34968 && 
b[34969] == 34969 && 
b[34970] == 34970 && 
b[34971] == 34971 && 
b[34972] == 34972 && 
b[34973] == 34973 && 
b[34974] == 34974 && 
b[34975] == 34975 && 
b[34976] == 34976 && 
b[34977] == 34977 && 
b[34978] == 34978 && 
b[34979] == 34979 && 
b[34980] == 34980 && 
b[34981] == 34981 && 
b[34982] == 34982 && 
b[34983] == 34983 && 
b[34984] == 34984 && 
b[34985] == 34985 && 
b[34986] == 34986 && 
b[34987] == 34987 && 
b[34988] == 34988 && 
b[34989] == 34989 && 
b[34990] == 34990 && 
b[34991] == 34991 && 
b[34992] == 34992 && 
b[34993] == 34993 && 
b[34994] == 34994 && 
b[34995] == 34995 && 
b[34996] == 34996 && 
b[34997] == 34997 && 
b[34998] == 34998 && 
b[34999] == 34999 && 
b[35000] == 35000 && 
b[35001] == 35001 && 
b[35002] == 35002 && 
b[35003] == 35003 && 
b[35004] == 35004 && 
b[35005] == 35005 && 
b[35006] == 35006 && 
b[35007] == 35007 && 
b[35008] == 35008 && 
b[35009] == 35009 && 
b[35010] == 35010 && 
b[35011] == 35011 && 
b[35012] == 35012 && 
b[35013] == 35013 && 
b[35014] == 35014 && 
b[35015] == 35015 && 
b[35016] == 35016 && 
b[35017] == 35017 && 
b[35018] == 35018 && 
b[35019] == 35019 && 
b[35020] == 35020 && 
b[35021] == 35021 && 
b[35022] == 35022 && 
b[35023] == 35023 && 
b[35024] == 35024 && 
b[35025] == 35025 && 
b[35026] == 35026 && 
b[35027] == 35027 && 
b[35028] == 35028 && 
b[35029] == 35029 && 
b[35030] == 35030 && 
b[35031] == 35031 && 
b[35032] == 35032 && 
b[35033] == 35033 && 
b[35034] == 35034 && 
b[35035] == 35035 && 
b[35036] == 35036 && 
b[35037] == 35037 && 
b[35038] == 35038 && 
b[35039] == 35039 && 
b[35040] == 35040 && 
b[35041] == 35041 && 
b[35042] == 35042 && 
b[35043] == 35043 && 
b[35044] == 35044 && 
b[35045] == 35045 && 
b[35046] == 35046 && 
b[35047] == 35047 && 
b[35048] == 35048 && 
b[35049] == 35049 && 
b[35050] == 35050 && 
b[35051] == 35051 && 
b[35052] == 35052 && 
b[35053] == 35053 && 
b[35054] == 35054 && 
b[35055] == 35055 && 
b[35056] == 35056 && 
b[35057] == 35057 && 
b[35058] == 35058 && 
b[35059] == 35059 && 
b[35060] == 35060 && 
b[35061] == 35061 && 
b[35062] == 35062 && 
b[35063] == 35063 && 
b[35064] == 35064 && 
b[35065] == 35065 && 
b[35066] == 35066 && 
b[35067] == 35067 && 
b[35068] == 35068 && 
b[35069] == 35069 && 
b[35070] == 35070 && 
b[35071] == 35071 && 
b[35072] == 35072 && 
b[35073] == 35073 && 
b[35074] == 35074 && 
b[35075] == 35075 && 
b[35076] == 35076 && 
b[35077] == 35077 && 
b[35078] == 35078 && 
b[35079] == 35079 && 
b[35080] == 35080 && 
b[35081] == 35081 && 
b[35082] == 35082 && 
b[35083] == 35083 && 
b[35084] == 35084 && 
b[35085] == 35085 && 
b[35086] == 35086 && 
b[35087] == 35087 && 
b[35088] == 35088 && 
b[35089] == 35089 && 
b[35090] == 35090 && 
b[35091] == 35091 && 
b[35092] == 35092 && 
b[35093] == 35093 && 
b[35094] == 35094 && 
b[35095] == 35095 && 
b[35096] == 35096 && 
b[35097] == 35097 && 
b[35098] == 35098 && 
b[35099] == 35099 && 
b[35100] == 35100 && 
b[35101] == 35101 && 
b[35102] == 35102 && 
b[35103] == 35103 && 
b[35104] == 35104 && 
b[35105] == 35105 && 
b[35106] == 35106 && 
b[35107] == 35107 && 
b[35108] == 35108 && 
b[35109] == 35109 && 
b[35110] == 35110 && 
b[35111] == 35111 && 
b[35112] == 35112 && 
b[35113] == 35113 && 
b[35114] == 35114 && 
b[35115] == 35115 && 
b[35116] == 35116 && 
b[35117] == 35117 && 
b[35118] == 35118 && 
b[35119] == 35119 && 
b[35120] == 35120 && 
b[35121] == 35121 && 
b[35122] == 35122 && 
b[35123] == 35123 && 
b[35124] == 35124 && 
b[35125] == 35125 && 
b[35126] == 35126 && 
b[35127] == 35127 && 
b[35128] == 35128 && 
b[35129] == 35129 && 
b[35130] == 35130 && 
b[35131] == 35131 && 
b[35132] == 35132 && 
b[35133] == 35133 && 
b[35134] == 35134 && 
b[35135] == 35135 && 
b[35136] == 35136 && 
b[35137] == 35137 && 
b[35138] == 35138 && 
b[35139] == 35139 && 
b[35140] == 35140 && 
b[35141] == 35141 && 
b[35142] == 35142 && 
b[35143] == 35143 && 
b[35144] == 35144 && 
b[35145] == 35145 && 
b[35146] == 35146 && 
b[35147] == 35147 && 
b[35148] == 35148 && 
b[35149] == 35149 && 
b[35150] == 35150 && 
b[35151] == 35151 && 
b[35152] == 35152 && 
b[35153] == 35153 && 
b[35154] == 35154 && 
b[35155] == 35155 && 
b[35156] == 35156 && 
b[35157] == 35157 && 
b[35158] == 35158 && 
b[35159] == 35159 && 
b[35160] == 35160 && 
b[35161] == 35161 && 
b[35162] == 35162 && 
b[35163] == 35163 && 
b[35164] == 35164 && 
b[35165] == 35165 && 
b[35166] == 35166 && 
b[35167] == 35167 && 
b[35168] == 35168 && 
b[35169] == 35169 && 
b[35170] == 35170 && 
b[35171] == 35171 && 
b[35172] == 35172 && 
b[35173] == 35173 && 
b[35174] == 35174 && 
b[35175] == 35175 && 
b[35176] == 35176 && 
b[35177] == 35177 && 
b[35178] == 35178 && 
b[35179] == 35179 && 
b[35180] == 35180 && 
b[35181] == 35181 && 
b[35182] == 35182 && 
b[35183] == 35183 && 
b[35184] == 35184 && 
b[35185] == 35185 && 
b[35186] == 35186 && 
b[35187] == 35187 && 
b[35188] == 35188 && 
b[35189] == 35189 && 
b[35190] == 35190 && 
b[35191] == 35191 && 
b[35192] == 35192 && 
b[35193] == 35193 && 
b[35194] == 35194 && 
b[35195] == 35195 && 
b[35196] == 35196 && 
b[35197] == 35197 && 
b[35198] == 35198 && 
b[35199] == 35199 && 
b[35200] == 35200 && 
b[35201] == 35201 && 
b[35202] == 35202 && 
b[35203] == 35203 && 
b[35204] == 35204 && 
b[35205] == 35205 && 
b[35206] == 35206 && 
b[35207] == 35207 && 
b[35208] == 35208 && 
b[35209] == 35209 && 
b[35210] == 35210 && 
b[35211] == 35211 && 
b[35212] == 35212 && 
b[35213] == 35213 && 
b[35214] == 35214 && 
b[35215] == 35215 && 
b[35216] == 35216 && 
b[35217] == 35217 && 
b[35218] == 35218 && 
b[35219] == 35219 && 
b[35220] == 35220 && 
b[35221] == 35221 && 
b[35222] == 35222 && 
b[35223] == 35223 && 
b[35224] == 35224 && 
b[35225] == 35225 && 
b[35226] == 35226 && 
b[35227] == 35227 && 
b[35228] == 35228 && 
b[35229] == 35229 && 
b[35230] == 35230 && 
b[35231] == 35231 && 
b[35232] == 35232 && 
b[35233] == 35233 && 
b[35234] == 35234 && 
b[35235] == 35235 && 
b[35236] == 35236 && 
b[35237] == 35237 && 
b[35238] == 35238 && 
b[35239] == 35239 && 
b[35240] == 35240 && 
b[35241] == 35241 && 
b[35242] == 35242 && 
b[35243] == 35243 && 
b[35244] == 35244 && 
b[35245] == 35245 && 
b[35246] == 35246 && 
b[35247] == 35247 && 
b[35248] == 35248 && 
b[35249] == 35249 && 
b[35250] == 35250 && 
b[35251] == 35251 && 
b[35252] == 35252 && 
b[35253] == 35253 && 
b[35254] == 35254 && 
b[35255] == 35255 && 
b[35256] == 35256 && 
b[35257] == 35257 && 
b[35258] == 35258 && 
b[35259] == 35259 && 
b[35260] == 35260 && 
b[35261] == 35261 && 
b[35262] == 35262 && 
b[35263] == 35263 && 
b[35264] == 35264 && 
b[35265] == 35265 && 
b[35266] == 35266 && 
b[35267] == 35267 && 
b[35268] == 35268 && 
b[35269] == 35269 && 
b[35270] == 35270 && 
b[35271] == 35271 && 
b[35272] == 35272 && 
b[35273] == 35273 && 
b[35274] == 35274 && 
b[35275] == 35275 && 
b[35276] == 35276 && 
b[35277] == 35277 && 
b[35278] == 35278 && 
b[35279] == 35279 && 
b[35280] == 35280 && 
b[35281] == 35281 && 
b[35282] == 35282 && 
b[35283] == 35283 && 
b[35284] == 35284 && 
b[35285] == 35285 && 
b[35286] == 35286 && 
b[35287] == 35287 && 
b[35288] == 35288 && 
b[35289] == 35289 && 
b[35290] == 35290 && 
b[35291] == 35291 && 
b[35292] == 35292 && 
b[35293] == 35293 && 
b[35294] == 35294 && 
b[35295] == 35295 && 
b[35296] == 35296 && 
b[35297] == 35297 && 
b[35298] == 35298 && 
b[35299] == 35299 && 
b[35300] == 35300 && 
b[35301] == 35301 && 
b[35302] == 35302 && 
b[35303] == 35303 && 
b[35304] == 35304 && 
b[35305] == 35305 && 
b[35306] == 35306 && 
b[35307] == 35307 && 
b[35308] == 35308 && 
b[35309] == 35309 && 
b[35310] == 35310 && 
b[35311] == 35311 && 
b[35312] == 35312 && 
b[35313] == 35313 && 
b[35314] == 35314 && 
b[35315] == 35315 && 
b[35316] == 35316 && 
b[35317] == 35317 && 
b[35318] == 35318 && 
b[35319] == 35319 && 
b[35320] == 35320 && 
b[35321] == 35321 && 
b[35322] == 35322 && 
b[35323] == 35323 && 
b[35324] == 35324 && 
b[35325] == 35325 && 
b[35326] == 35326 && 
b[35327] == 35327 && 
b[35328] == 35328 && 
b[35329] == 35329 && 
b[35330] == 35330 && 
b[35331] == 35331 && 
b[35332] == 35332 && 
b[35333] == 35333 && 
b[35334] == 35334 && 
b[35335] == 35335 && 
b[35336] == 35336 && 
b[35337] == 35337 && 
b[35338] == 35338 && 
b[35339] == 35339 && 
b[35340] == 35340 && 
b[35341] == 35341 && 
b[35342] == 35342 && 
b[35343] == 35343 && 
b[35344] == 35344 && 
b[35345] == 35345 && 
b[35346] == 35346 && 
b[35347] == 35347 && 
b[35348] == 35348 && 
b[35349] == 35349 && 
b[35350] == 35350 && 
b[35351] == 35351 && 
b[35352] == 35352 && 
b[35353] == 35353 && 
b[35354] == 35354 && 
b[35355] == 35355 && 
b[35356] == 35356 && 
b[35357] == 35357 && 
b[35358] == 35358 && 
b[35359] == 35359 && 
b[35360] == 35360 && 
b[35361] == 35361 && 
b[35362] == 35362 && 
b[35363] == 35363 && 
b[35364] == 35364 && 
b[35365] == 35365 && 
b[35366] == 35366 && 
b[35367] == 35367 && 
b[35368] == 35368 && 
b[35369] == 35369 && 
b[35370] == 35370 && 
b[35371] == 35371 && 
b[35372] == 35372 && 
b[35373] == 35373 && 
b[35374] == 35374 && 
b[35375] == 35375 && 
b[35376] == 35376 && 
b[35377] == 35377 && 
b[35378] == 35378 && 
b[35379] == 35379 && 
b[35380] == 35380 && 
b[35381] == 35381 && 
b[35382] == 35382 && 
b[35383] == 35383 && 
b[35384] == 35384 && 
b[35385] == 35385 && 
b[35386] == 35386 && 
b[35387] == 35387 && 
b[35388] == 35388 && 
b[35389] == 35389 && 
b[35390] == 35390 && 
b[35391] == 35391 && 
b[35392] == 35392 && 
b[35393] == 35393 && 
b[35394] == 35394 && 
b[35395] == 35395 && 
b[35396] == 35396 && 
b[35397] == 35397 && 
b[35398] == 35398 && 
b[35399] == 35399 && 
b[35400] == 35400 && 
b[35401] == 35401 && 
b[35402] == 35402 && 
b[35403] == 35403 && 
b[35404] == 35404 && 
b[35405] == 35405 && 
b[35406] == 35406 && 
b[35407] == 35407 && 
b[35408] == 35408 && 
b[35409] == 35409 && 
b[35410] == 35410 && 
b[35411] == 35411 && 
b[35412] == 35412 && 
b[35413] == 35413 && 
b[35414] == 35414 && 
b[35415] == 35415 && 
b[35416] == 35416 && 
b[35417] == 35417 && 
b[35418] == 35418 && 
b[35419] == 35419 && 
b[35420] == 35420 && 
b[35421] == 35421 && 
b[35422] == 35422 && 
b[35423] == 35423 && 
b[35424] == 35424 && 
b[35425] == 35425 && 
b[35426] == 35426 && 
b[35427] == 35427 && 
b[35428] == 35428 && 
b[35429] == 35429 && 
b[35430] == 35430 && 
b[35431] == 35431 && 
b[35432] == 35432 && 
b[35433] == 35433 && 
b[35434] == 35434 && 
b[35435] == 35435 && 
b[35436] == 35436 && 
b[35437] == 35437 && 
b[35438] == 35438 && 
b[35439] == 35439 && 
b[35440] == 35440 && 
b[35441] == 35441 && 
b[35442] == 35442 && 
b[35443] == 35443 && 
b[35444] == 35444 && 
b[35445] == 35445 && 
b[35446] == 35446 && 
b[35447] == 35447 && 
b[35448] == 35448 && 
b[35449] == 35449 && 
b[35450] == 35450 && 
b[35451] == 35451 && 
b[35452] == 35452 && 
b[35453] == 35453 && 
b[35454] == 35454 && 
b[35455] == 35455 && 
b[35456] == 35456 && 
b[35457] == 35457 && 
b[35458] == 35458 && 
b[35459] == 35459 && 
b[35460] == 35460 && 
b[35461] == 35461 && 
b[35462] == 35462 && 
b[35463] == 35463 && 
b[35464] == 35464 && 
b[35465] == 35465 && 
b[35466] == 35466 && 
b[35467] == 35467 && 
b[35468] == 35468 && 
b[35469] == 35469 && 
b[35470] == 35470 && 
b[35471] == 35471 && 
b[35472] == 35472 && 
b[35473] == 35473 && 
b[35474] == 35474 && 
b[35475] == 35475 && 
b[35476] == 35476 && 
b[35477] == 35477 && 
b[35478] == 35478 && 
b[35479] == 35479 && 
b[35480] == 35480 && 
b[35481] == 35481 && 
b[35482] == 35482 && 
b[35483] == 35483 && 
b[35484] == 35484 && 
b[35485] == 35485 && 
b[35486] == 35486 && 
b[35487] == 35487 && 
b[35488] == 35488 && 
b[35489] == 35489 && 
b[35490] == 35490 && 
b[35491] == 35491 && 
b[35492] == 35492 && 
b[35493] == 35493 && 
b[35494] == 35494 && 
b[35495] == 35495 && 
b[35496] == 35496 && 
b[35497] == 35497 && 
b[35498] == 35498 && 
b[35499] == 35499 && 
b[35500] == 35500 && 
b[35501] == 35501 && 
b[35502] == 35502 && 
b[35503] == 35503 && 
b[35504] == 35504 && 
b[35505] == 35505 && 
b[35506] == 35506 && 
b[35507] == 35507 && 
b[35508] == 35508 && 
b[35509] == 35509 && 
b[35510] == 35510 && 
b[35511] == 35511 && 
b[35512] == 35512 && 
b[35513] == 35513 && 
b[35514] == 35514 && 
b[35515] == 35515 && 
b[35516] == 35516 && 
b[35517] == 35517 && 
b[35518] == 35518 && 
b[35519] == 35519 && 
b[35520] == 35520 && 
b[35521] == 35521 && 
b[35522] == 35522 && 
b[35523] == 35523 && 
b[35524] == 35524 && 
b[35525] == 35525 && 
b[35526] == 35526 && 
b[35527] == 35527 && 
b[35528] == 35528 && 
b[35529] == 35529 && 
b[35530] == 35530 && 
b[35531] == 35531 && 
b[35532] == 35532 && 
b[35533] == 35533 && 
b[35534] == 35534 && 
b[35535] == 35535 && 
b[35536] == 35536 && 
b[35537] == 35537 && 
b[35538] == 35538 && 
b[35539] == 35539 && 
b[35540] == 35540 && 
b[35541] == 35541 && 
b[35542] == 35542 && 
b[35543] == 35543 && 
b[35544] == 35544 && 
b[35545] == 35545 && 
b[35546] == 35546 && 
b[35547] == 35547 && 
b[35548] == 35548 && 
b[35549] == 35549 && 
b[35550] == 35550 && 
b[35551] == 35551 && 
b[35552] == 35552 && 
b[35553] == 35553 && 
b[35554] == 35554 && 
b[35555] == 35555 && 
b[35556] == 35556 && 
b[35557] == 35557 && 
b[35558] == 35558 && 
b[35559] == 35559 && 
b[35560] == 35560 && 
b[35561] == 35561 && 
b[35562] == 35562 && 
b[35563] == 35563 && 
b[35564] == 35564 && 
b[35565] == 35565 && 
b[35566] == 35566 && 
b[35567] == 35567 && 
b[35568] == 35568 && 
b[35569] == 35569 && 
b[35570] == 35570 && 
b[35571] == 35571 && 
b[35572] == 35572 && 
b[35573] == 35573 && 
b[35574] == 35574 && 
b[35575] == 35575 && 
b[35576] == 35576 && 
b[35577] == 35577 && 
b[35578] == 35578 && 
b[35579] == 35579 && 
b[35580] == 35580 && 
b[35581] == 35581 && 
b[35582] == 35582 && 
b[35583] == 35583 && 
b[35584] == 35584 && 
b[35585] == 35585 && 
b[35586] == 35586 && 
b[35587] == 35587 && 
b[35588] == 35588 && 
b[35589] == 35589 && 
b[35590] == 35590 && 
b[35591] == 35591 && 
b[35592] == 35592 && 
b[35593] == 35593 && 
b[35594] == 35594 && 
b[35595] == 35595 && 
b[35596] == 35596 && 
b[35597] == 35597 && 
b[35598] == 35598 && 
b[35599] == 35599 && 
b[35600] == 35600 && 
b[35601] == 35601 && 
b[35602] == 35602 && 
b[35603] == 35603 && 
b[35604] == 35604 && 
b[35605] == 35605 && 
b[35606] == 35606 && 
b[35607] == 35607 && 
b[35608] == 35608 && 
b[35609] == 35609 && 
b[35610] == 35610 && 
b[35611] == 35611 && 
b[35612] == 35612 && 
b[35613] == 35613 && 
b[35614] == 35614 && 
b[35615] == 35615 && 
b[35616] == 35616 && 
b[35617] == 35617 && 
b[35618] == 35618 && 
b[35619] == 35619 && 
b[35620] == 35620 && 
b[35621] == 35621 && 
b[35622] == 35622 && 
b[35623] == 35623 && 
b[35624] == 35624 && 
b[35625] == 35625 && 
b[35626] == 35626 && 
b[35627] == 35627 && 
b[35628] == 35628 && 
b[35629] == 35629 && 
b[35630] == 35630 && 
b[35631] == 35631 && 
b[35632] == 35632 && 
b[35633] == 35633 && 
b[35634] == 35634 && 
b[35635] == 35635 && 
b[35636] == 35636 && 
b[35637] == 35637 && 
b[35638] == 35638 && 
b[35639] == 35639 && 
b[35640] == 35640 && 
b[35641] == 35641 && 
b[35642] == 35642 && 
b[35643] == 35643 && 
b[35644] == 35644 && 
b[35645] == 35645 && 
b[35646] == 35646 && 
b[35647] == 35647 && 
b[35648] == 35648 && 
b[35649] == 35649 && 
b[35650] == 35650 && 
b[35651] == 35651 && 
b[35652] == 35652 && 
b[35653] == 35653 && 
b[35654] == 35654 && 
b[35655] == 35655 && 
b[35656] == 35656 && 
b[35657] == 35657 && 
b[35658] == 35658 && 
b[35659] == 35659 && 
b[35660] == 35660 && 
b[35661] == 35661 && 
b[35662] == 35662 && 
b[35663] == 35663 && 
b[35664] == 35664 && 
b[35665] == 35665 && 
b[35666] == 35666 && 
b[35667] == 35667 && 
b[35668] == 35668 && 
b[35669] == 35669 && 
b[35670] == 35670 && 
b[35671] == 35671 && 
b[35672] == 35672 && 
b[35673] == 35673 && 
b[35674] == 35674 && 
b[35675] == 35675 && 
b[35676] == 35676 && 
b[35677] == 35677 && 
b[35678] == 35678 && 
b[35679] == 35679 && 
b[35680] == 35680 && 
b[35681] == 35681 && 
b[35682] == 35682 && 
b[35683] == 35683 && 
b[35684] == 35684 && 
b[35685] == 35685 && 
b[35686] == 35686 && 
b[35687] == 35687 && 
b[35688] == 35688 && 
b[35689] == 35689 && 
b[35690] == 35690 && 
b[35691] == 35691 && 
b[35692] == 35692 && 
b[35693] == 35693 && 
b[35694] == 35694 && 
b[35695] == 35695 && 
b[35696] == 35696 && 
b[35697] == 35697 && 
b[35698] == 35698 && 
b[35699] == 35699 && 
b[35700] == 35700 && 
b[35701] == 35701 && 
b[35702] == 35702 && 
b[35703] == 35703 && 
b[35704] == 35704 && 
b[35705] == 35705 && 
b[35706] == 35706 && 
b[35707] == 35707 && 
b[35708] == 35708 && 
b[35709] == 35709 && 
b[35710] == 35710 && 
b[35711] == 35711 && 
b[35712] == 35712 && 
b[35713] == 35713 && 
b[35714] == 35714 && 
b[35715] == 35715 && 
b[35716] == 35716 && 
b[35717] == 35717 && 
b[35718] == 35718 && 
b[35719] == 35719 && 
b[35720] == 35720 && 
b[35721] == 35721 && 
b[35722] == 35722 && 
b[35723] == 35723 && 
b[35724] == 35724 && 
b[35725] == 35725 && 
b[35726] == 35726 && 
b[35727] == 35727 && 
b[35728] == 35728 && 
b[35729] == 35729 && 
b[35730] == 35730 && 
b[35731] == 35731 && 
b[35732] == 35732 && 
b[35733] == 35733 && 
b[35734] == 35734 && 
b[35735] == 35735 && 
b[35736] == 35736 && 
b[35737] == 35737 && 
b[35738] == 35738 && 
b[35739] == 35739 && 
b[35740] == 35740 && 
b[35741] == 35741 && 
b[35742] == 35742 && 
b[35743] == 35743 && 
b[35744] == 35744 && 
b[35745] == 35745 && 
b[35746] == 35746 && 
b[35747] == 35747 && 
b[35748] == 35748 && 
b[35749] == 35749 && 
b[35750] == 35750 && 
b[35751] == 35751 && 
b[35752] == 35752 && 
b[35753] == 35753 && 
b[35754] == 35754 && 
b[35755] == 35755 && 
b[35756] == 35756 && 
b[35757] == 35757 && 
b[35758] == 35758 && 
b[35759] == 35759 && 
b[35760] == 35760 && 
b[35761] == 35761 && 
b[35762] == 35762 && 
b[35763] == 35763 && 
b[35764] == 35764 && 
b[35765] == 35765 && 
b[35766] == 35766 && 
b[35767] == 35767 && 
b[35768] == 35768 && 
b[35769] == 35769 && 
b[35770] == 35770 && 
b[35771] == 35771 && 
b[35772] == 35772 && 
b[35773] == 35773 && 
b[35774] == 35774 && 
b[35775] == 35775 && 
b[35776] == 35776 && 
b[35777] == 35777 && 
b[35778] == 35778 && 
b[35779] == 35779 && 
b[35780] == 35780 && 
b[35781] == 35781 && 
b[35782] == 35782 && 
b[35783] == 35783 && 
b[35784] == 35784 && 
b[35785] == 35785 && 
b[35786] == 35786 && 
b[35787] == 35787 && 
b[35788] == 35788 && 
b[35789] == 35789 && 
b[35790] == 35790 && 
b[35791] == 35791 && 
b[35792] == 35792 && 
b[35793] == 35793 && 
b[35794] == 35794 && 
b[35795] == 35795 && 
b[35796] == 35796 && 
b[35797] == 35797 && 
b[35798] == 35798 && 
b[35799] == 35799 && 
b[35800] == 35800 && 
b[35801] == 35801 && 
b[35802] == 35802 && 
b[35803] == 35803 && 
b[35804] == 35804 && 
b[35805] == 35805 && 
b[35806] == 35806 && 
b[35807] == 35807 && 
b[35808] == 35808 && 
b[35809] == 35809 && 
b[35810] == 35810 && 
b[35811] == 35811 && 
b[35812] == 35812 && 
b[35813] == 35813 && 
b[35814] == 35814 && 
b[35815] == 35815 && 
b[35816] == 35816 && 
b[35817] == 35817 && 
b[35818] == 35818 && 
b[35819] == 35819 && 
b[35820] == 35820 && 
b[35821] == 35821 && 
b[35822] == 35822 && 
b[35823] == 35823 && 
b[35824] == 35824 && 
b[35825] == 35825 && 
b[35826] == 35826 && 
b[35827] == 35827 && 
b[35828] == 35828 && 
b[35829] == 35829 && 
b[35830] == 35830 && 
b[35831] == 35831 && 
b[35832] == 35832 && 
b[35833] == 35833 && 
b[35834] == 35834 && 
b[35835] == 35835 && 
b[35836] == 35836 && 
b[35837] == 35837 && 
b[35838] == 35838 && 
b[35839] == 35839 && 
b[35840] == 35840 && 
b[35841] == 35841 && 
b[35842] == 35842 && 
b[35843] == 35843 && 
b[35844] == 35844 && 
b[35845] == 35845 && 
b[35846] == 35846 && 
b[35847] == 35847 && 
b[35848] == 35848 && 
b[35849] == 35849 && 
b[35850] == 35850 && 
b[35851] == 35851 && 
b[35852] == 35852 && 
b[35853] == 35853 && 
b[35854] == 35854 && 
b[35855] == 35855 && 
b[35856] == 35856 && 
b[35857] == 35857 && 
b[35858] == 35858 && 
b[35859] == 35859 && 
b[35860] == 35860 && 
b[35861] == 35861 && 
b[35862] == 35862 && 
b[35863] == 35863 && 
b[35864] == 35864 && 
b[35865] == 35865 && 
b[35866] == 35866 && 
b[35867] == 35867 && 
b[35868] == 35868 && 
b[35869] == 35869 && 
b[35870] == 35870 && 
b[35871] == 35871 && 
b[35872] == 35872 && 
b[35873] == 35873 && 
b[35874] == 35874 && 
b[35875] == 35875 && 
b[35876] == 35876 && 
b[35877] == 35877 && 
b[35878] == 35878 && 
b[35879] == 35879 && 
b[35880] == 35880 && 
b[35881] == 35881 && 
b[35882] == 35882 && 
b[35883] == 35883 && 
b[35884] == 35884 && 
b[35885] == 35885 && 
b[35886] == 35886 && 
b[35887] == 35887 && 
b[35888] == 35888 && 
b[35889] == 35889 && 
b[35890] == 35890 && 
b[35891] == 35891 && 
b[35892] == 35892 && 
b[35893] == 35893 && 
b[35894] == 35894 && 
b[35895] == 35895 && 
b[35896] == 35896 && 
b[35897] == 35897 && 
b[35898] == 35898 && 
b[35899] == 35899 && 
b[35900] == 35900 && 
b[35901] == 35901 && 
b[35902] == 35902 && 
b[35903] == 35903 && 
b[35904] == 35904 && 
b[35905] == 35905 && 
b[35906] == 35906 && 
b[35907] == 35907 && 
b[35908] == 35908 && 
b[35909] == 35909 && 
b[35910] == 35910 && 
b[35911] == 35911 && 
b[35912] == 35912 && 
b[35913] == 35913 && 
b[35914] == 35914 && 
b[35915] == 35915 && 
b[35916] == 35916 && 
b[35917] == 35917 && 
b[35918] == 35918 && 
b[35919] == 35919 && 
b[35920] == 35920 && 
b[35921] == 35921 && 
b[35922] == 35922 && 
b[35923] == 35923 && 
b[35924] == 35924 && 
b[35925] == 35925 && 
b[35926] == 35926 && 
b[35927] == 35927 && 
b[35928] == 35928 && 
b[35929] == 35929 && 
b[35930] == 35930 && 
b[35931] == 35931 && 
b[35932] == 35932 && 
b[35933] == 35933 && 
b[35934] == 35934 && 
b[35935] == 35935 && 
b[35936] == 35936 && 
b[35937] == 35937 && 
b[35938] == 35938 && 
b[35939] == 35939 && 
b[35940] == 35940 && 
b[35941] == 35941 && 
b[35942] == 35942 && 
b[35943] == 35943 && 
b[35944] == 35944 && 
b[35945] == 35945 && 
b[35946] == 35946 && 
b[35947] == 35947 && 
b[35948] == 35948 && 
b[35949] == 35949 && 
b[35950] == 35950 && 
b[35951] == 35951 && 
b[35952] == 35952 && 
b[35953] == 35953 && 
b[35954] == 35954 && 
b[35955] == 35955 && 
b[35956] == 35956 && 
b[35957] == 35957 && 
b[35958] == 35958 && 
b[35959] == 35959 && 
b[35960] == 35960 && 
b[35961] == 35961 && 
b[35962] == 35962 && 
b[35963] == 35963 && 
b[35964] == 35964 && 
b[35965] == 35965 && 
b[35966] == 35966 && 
b[35967] == 35967 && 
b[35968] == 35968 && 
b[35969] == 35969 && 
b[35970] == 35970 && 
b[35971] == 35971 && 
b[35972] == 35972 && 
b[35973] == 35973 && 
b[35974] == 35974 && 
b[35975] == 35975 && 
b[35976] == 35976 && 
b[35977] == 35977 && 
b[35978] == 35978 && 
b[35979] == 35979 && 
b[35980] == 35980 && 
b[35981] == 35981 && 
b[35982] == 35982 && 
b[35983] == 35983 && 
b[35984] == 35984 && 
b[35985] == 35985 && 
b[35986] == 35986 && 
b[35987] == 35987 && 
b[35988] == 35988 && 
b[35989] == 35989 && 
b[35990] == 35990 && 
b[35991] == 35991 && 
b[35992] == 35992 && 
b[35993] == 35993 && 
b[35994] == 35994 && 
b[35995] == 35995 && 
b[35996] == 35996 && 
b[35997] == 35997 && 
b[35998] == 35998 && 
b[35999] == 35999 && 
b[36000] == 36000 && 
b[36001] == 36001 && 
b[36002] == 36002 && 
b[36003] == 36003 && 
b[36004] == 36004 && 
b[36005] == 36005 && 
b[36006] == 36006 && 
b[36007] == 36007 && 
b[36008] == 36008 && 
b[36009] == 36009 && 
b[36010] == 36010 && 
b[36011] == 36011 && 
b[36012] == 36012 && 
b[36013] == 36013 && 
b[36014] == 36014 && 
b[36015] == 36015 && 
b[36016] == 36016 && 
b[36017] == 36017 && 
b[36018] == 36018 && 
b[36019] == 36019 && 
b[36020] == 36020 && 
b[36021] == 36021 && 
b[36022] == 36022 && 
b[36023] == 36023 && 
b[36024] == 36024 && 
b[36025] == 36025 && 
b[36026] == 36026 && 
b[36027] == 36027 && 
b[36028] == 36028 && 
b[36029] == 36029 && 
b[36030] == 36030 && 
b[36031] == 36031 && 
b[36032] == 36032 && 
b[36033] == 36033 && 
b[36034] == 36034 && 
b[36035] == 36035 && 
b[36036] == 36036 && 
b[36037] == 36037 && 
b[36038] == 36038 && 
b[36039] == 36039 && 
b[36040] == 36040 && 
b[36041] == 36041 && 
b[36042] == 36042 && 
b[36043] == 36043 && 
b[36044] == 36044 && 
b[36045] == 36045 && 
b[36046] == 36046 && 
b[36047] == 36047 && 
b[36048] == 36048 && 
b[36049] == 36049 && 
b[36050] == 36050 && 
b[36051] == 36051 && 
b[36052] == 36052 && 
b[36053] == 36053 && 
b[36054] == 36054 && 
b[36055] == 36055 && 
b[36056] == 36056 && 
b[36057] == 36057 && 
b[36058] == 36058 && 
b[36059] == 36059 && 
b[36060] == 36060 && 
b[36061] == 36061 && 
b[36062] == 36062 && 
b[36063] == 36063 && 
b[36064] == 36064 && 
b[36065] == 36065 && 
b[36066] == 36066 && 
b[36067] == 36067 && 
b[36068] == 36068 && 
b[36069] == 36069 && 
b[36070] == 36070 && 
b[36071] == 36071 && 
b[36072] == 36072 && 
b[36073] == 36073 && 
b[36074] == 36074 && 
b[36075] == 36075 && 
b[36076] == 36076 && 
b[36077] == 36077 && 
b[36078] == 36078 && 
b[36079] == 36079 && 
b[36080] == 36080 && 
b[36081] == 36081 && 
b[36082] == 36082 && 
b[36083] == 36083 && 
b[36084] == 36084 && 
b[36085] == 36085 && 
b[36086] == 36086 && 
b[36087] == 36087 && 
b[36088] == 36088 && 
b[36089] == 36089 && 
b[36090] == 36090 && 
b[36091] == 36091 && 
b[36092] == 36092 && 
b[36093] == 36093 && 
b[36094] == 36094 && 
b[36095] == 36095 && 
b[36096] == 36096 && 
b[36097] == 36097 && 
b[36098] == 36098 && 
b[36099] == 36099 && 
b[36100] == 36100 && 
b[36101] == 36101 && 
b[36102] == 36102 && 
b[36103] == 36103 && 
b[36104] == 36104 && 
b[36105] == 36105 && 
b[36106] == 36106 && 
b[36107] == 36107 && 
b[36108] == 36108 && 
b[36109] == 36109 && 
b[36110] == 36110 && 
b[36111] == 36111 && 
b[36112] == 36112 && 
b[36113] == 36113 && 
b[36114] == 36114 && 
b[36115] == 36115 && 
b[36116] == 36116 && 
b[36117] == 36117 && 
b[36118] == 36118 && 
b[36119] == 36119 && 
b[36120] == 36120 && 
b[36121] == 36121 && 
b[36122] == 36122 && 
b[36123] == 36123 && 
b[36124] == 36124 && 
b[36125] == 36125 && 
b[36126] == 36126 && 
b[36127] == 36127 && 
b[36128] == 36128 && 
b[36129] == 36129 && 
b[36130] == 36130 && 
b[36131] == 36131 && 
b[36132] == 36132 && 
b[36133] == 36133 && 
b[36134] == 36134 && 
b[36135] == 36135 && 
b[36136] == 36136 && 
b[36137] == 36137 && 
b[36138] == 36138 && 
b[36139] == 36139 && 
b[36140] == 36140 && 
b[36141] == 36141 && 
b[36142] == 36142 && 
b[36143] == 36143 && 
b[36144] == 36144 && 
b[36145] == 36145 && 
b[36146] == 36146 && 
b[36147] == 36147 && 
b[36148] == 36148 && 
b[36149] == 36149 && 
b[36150] == 36150 && 
b[36151] == 36151 && 
b[36152] == 36152 && 
b[36153] == 36153 && 
b[36154] == 36154 && 
b[36155] == 36155 && 
b[36156] == 36156 && 
b[36157] == 36157 && 
b[36158] == 36158 && 
b[36159] == 36159 && 
b[36160] == 36160 && 
b[36161] == 36161 && 
b[36162] == 36162 && 
b[36163] == 36163 && 
b[36164] == 36164 && 
b[36165] == 36165 && 
b[36166] == 36166 && 
b[36167] == 36167 && 
b[36168] == 36168 && 
b[36169] == 36169 && 
b[36170] == 36170 && 
b[36171] == 36171 && 
b[36172] == 36172 && 
b[36173] == 36173 && 
b[36174] == 36174 && 
b[36175] == 36175 && 
b[36176] == 36176 && 
b[36177] == 36177 && 
b[36178] == 36178 && 
b[36179] == 36179 && 
b[36180] == 36180 && 
b[36181] == 36181 && 
b[36182] == 36182 && 
b[36183] == 36183 && 
b[36184] == 36184 && 
b[36185] == 36185 && 
b[36186] == 36186 && 
b[36187] == 36187 && 
b[36188] == 36188 && 
b[36189] == 36189 && 
b[36190] == 36190 && 
b[36191] == 36191 && 
b[36192] == 36192 && 
b[36193] == 36193 && 
b[36194] == 36194 && 
b[36195] == 36195 && 
b[36196] == 36196 && 
b[36197] == 36197 && 
b[36198] == 36198 && 
b[36199] == 36199 && 
b[36200] == 36200 && 
b[36201] == 36201 && 
b[36202] == 36202 && 
b[36203] == 36203 && 
b[36204] == 36204 && 
b[36205] == 36205 && 
b[36206] == 36206 && 
b[36207] == 36207 && 
b[36208] == 36208 && 
b[36209] == 36209 && 
b[36210] == 36210 && 
b[36211] == 36211 && 
b[36212] == 36212 && 
b[36213] == 36213 && 
b[36214] == 36214 && 
b[36215] == 36215 && 
b[36216] == 36216 && 
b[36217] == 36217 && 
b[36218] == 36218 && 
b[36219] == 36219 && 
b[36220] == 36220 && 
b[36221] == 36221 && 
b[36222] == 36222 && 
b[36223] == 36223 && 
b[36224] == 36224 && 
b[36225] == 36225 && 
b[36226] == 36226 && 
b[36227] == 36227 && 
b[36228] == 36228 && 
b[36229] == 36229 && 
b[36230] == 36230 && 
b[36231] == 36231 && 
b[36232] == 36232 && 
b[36233] == 36233 && 
b[36234] == 36234 && 
b[36235] == 36235 && 
b[36236] == 36236 && 
b[36237] == 36237 && 
b[36238] == 36238 && 
b[36239] == 36239 && 
b[36240] == 36240 && 
b[36241] == 36241 && 
b[36242] == 36242 && 
b[36243] == 36243 && 
b[36244] == 36244 && 
b[36245] == 36245 && 
b[36246] == 36246 && 
b[36247] == 36247 && 
b[36248] == 36248 && 
b[36249] == 36249 && 
b[36250] == 36250 && 
b[36251] == 36251 && 
b[36252] == 36252 && 
b[36253] == 36253 && 
b[36254] == 36254 && 
b[36255] == 36255 && 
b[36256] == 36256 && 
b[36257] == 36257 && 
b[36258] == 36258 && 
b[36259] == 36259 && 
b[36260] == 36260 && 
b[36261] == 36261 && 
b[36262] == 36262 && 
b[36263] == 36263 && 
b[36264] == 36264 && 
b[36265] == 36265 && 
b[36266] == 36266 && 
b[36267] == 36267 && 
b[36268] == 36268 && 
b[36269] == 36269 && 
b[36270] == 36270 && 
b[36271] == 36271 && 
b[36272] == 36272 && 
b[36273] == 36273 && 
b[36274] == 36274 && 
b[36275] == 36275 && 
b[36276] == 36276 && 
b[36277] == 36277 && 
b[36278] == 36278 && 
b[36279] == 36279 && 
b[36280] == 36280 && 
b[36281] == 36281 && 
b[36282] == 36282 && 
b[36283] == 36283 && 
b[36284] == 36284 && 
b[36285] == 36285 && 
b[36286] == 36286 && 
b[36287] == 36287 && 
b[36288] == 36288 && 
b[36289] == 36289 && 
b[36290] == 36290 && 
b[36291] == 36291 && 
b[36292] == 36292 && 
b[36293] == 36293 && 
b[36294] == 36294 && 
b[36295] == 36295 && 
b[36296] == 36296 && 
b[36297] == 36297 && 
b[36298] == 36298 && 
b[36299] == 36299 && 
b[36300] == 36300 && 
b[36301] == 36301 && 
b[36302] == 36302 && 
b[36303] == 36303 && 
b[36304] == 36304 && 
b[36305] == 36305 && 
b[36306] == 36306 && 
b[36307] == 36307 && 
b[36308] == 36308 && 
b[36309] == 36309 && 
b[36310] == 36310 && 
b[36311] == 36311 && 
b[36312] == 36312 && 
b[36313] == 36313 && 
b[36314] == 36314 && 
b[36315] == 36315 && 
b[36316] == 36316 && 
b[36317] == 36317 && 
b[36318] == 36318 && 
b[36319] == 36319 && 
b[36320] == 36320 && 
b[36321] == 36321 && 
b[36322] == 36322 && 
b[36323] == 36323 && 
b[36324] == 36324 && 
b[36325] == 36325 && 
b[36326] == 36326 && 
b[36327] == 36327 && 
b[36328] == 36328 && 
b[36329] == 36329 && 
b[36330] == 36330 && 
b[36331] == 36331 && 
b[36332] == 36332 && 
b[36333] == 36333 && 
b[36334] == 36334 && 
b[36335] == 36335 && 
b[36336] == 36336 && 
b[36337] == 36337 && 
b[36338] == 36338 && 
b[36339] == 36339 && 
b[36340] == 36340 && 
b[36341] == 36341 && 
b[36342] == 36342 && 
b[36343] == 36343 && 
b[36344] == 36344 && 
b[36345] == 36345 && 
b[36346] == 36346 && 
b[36347] == 36347 && 
b[36348] == 36348 && 
b[36349] == 36349 && 
b[36350] == 36350 && 
b[36351] == 36351 && 
b[36352] == 36352 && 
b[36353] == 36353 && 
b[36354] == 36354 && 
b[36355] == 36355 && 
b[36356] == 36356 && 
b[36357] == 36357 && 
b[36358] == 36358 && 
b[36359] == 36359 && 
b[36360] == 36360 && 
b[36361] == 36361 && 
b[36362] == 36362 && 
b[36363] == 36363 && 
b[36364] == 36364 && 
b[36365] == 36365 && 
b[36366] == 36366 && 
b[36367] == 36367 && 
b[36368] == 36368 && 
b[36369] == 36369 && 
b[36370] == 36370 && 
b[36371] == 36371 && 
b[36372] == 36372 && 
b[36373] == 36373 && 
b[36374] == 36374 && 
b[36375] == 36375 && 
b[36376] == 36376 && 
b[36377] == 36377 && 
b[36378] == 36378 && 
b[36379] == 36379 && 
b[36380] == 36380 && 
b[36381] == 36381 && 
b[36382] == 36382 && 
b[36383] == 36383 && 
b[36384] == 36384 && 
b[36385] == 36385 && 
b[36386] == 36386 && 
b[36387] == 36387 && 
b[36388] == 36388 && 
b[36389] == 36389 && 
b[36390] == 36390 && 
b[36391] == 36391 && 
b[36392] == 36392 && 
b[36393] == 36393 && 
b[36394] == 36394 && 
b[36395] == 36395 && 
b[36396] == 36396 && 
b[36397] == 36397 && 
b[36398] == 36398 && 
b[36399] == 36399 && 
b[36400] == 36400 && 
b[36401] == 36401 && 
b[36402] == 36402 && 
b[36403] == 36403 && 
b[36404] == 36404 && 
b[36405] == 36405 && 
b[36406] == 36406 && 
b[36407] == 36407 && 
b[36408] == 36408 && 
b[36409] == 36409 && 
b[36410] == 36410 && 
b[36411] == 36411 && 
b[36412] == 36412 && 
b[36413] == 36413 && 
b[36414] == 36414 && 
b[36415] == 36415 && 
b[36416] == 36416 && 
b[36417] == 36417 && 
b[36418] == 36418 && 
b[36419] == 36419 && 
b[36420] == 36420 && 
b[36421] == 36421 && 
b[36422] == 36422 && 
b[36423] == 36423 && 
b[36424] == 36424 && 
b[36425] == 36425 && 
b[36426] == 36426 && 
b[36427] == 36427 && 
b[36428] == 36428 && 
b[36429] == 36429 && 
b[36430] == 36430 && 
b[36431] == 36431 && 
b[36432] == 36432 && 
b[36433] == 36433 && 
b[36434] == 36434 && 
b[36435] == 36435 && 
b[36436] == 36436 && 
b[36437] == 36437 && 
b[36438] == 36438 && 
b[36439] == 36439 && 
b[36440] == 36440 && 
b[36441] == 36441 && 
b[36442] == 36442 && 
b[36443] == 36443 && 
b[36444] == 36444 && 
b[36445] == 36445 && 
b[36446] == 36446 && 
b[36447] == 36447 && 
b[36448] == 36448 && 
b[36449] == 36449 && 
b[36450] == 36450 && 
b[36451] == 36451 && 
b[36452] == 36452 && 
b[36453] == 36453 && 
b[36454] == 36454 && 
b[36455] == 36455 && 
b[36456] == 36456 && 
b[36457] == 36457 && 
b[36458] == 36458 && 
b[36459] == 36459 && 
b[36460] == 36460 && 
b[36461] == 36461 && 
b[36462] == 36462 && 
b[36463] == 36463 && 
b[36464] == 36464 && 
b[36465] == 36465 && 
b[36466] == 36466 && 
b[36467] == 36467 && 
b[36468] == 36468 && 
b[36469] == 36469 && 
b[36470] == 36470 && 
b[36471] == 36471 && 
b[36472] == 36472 && 
b[36473] == 36473 && 
b[36474] == 36474 && 
b[36475] == 36475 && 
b[36476] == 36476 && 
b[36477] == 36477 && 
b[36478] == 36478 && 
b[36479] == 36479 && 
b[36480] == 36480 && 
b[36481] == 36481 && 
b[36482] == 36482 && 
b[36483] == 36483 && 
b[36484] == 36484 && 
b[36485] == 36485 && 
b[36486] == 36486 && 
b[36487] == 36487 && 
b[36488] == 36488 && 
b[36489] == 36489 && 
b[36490] == 36490 && 
b[36491] == 36491 && 
b[36492] == 36492 && 
b[36493] == 36493 && 
b[36494] == 36494 && 
b[36495] == 36495 && 
b[36496] == 36496 && 
b[36497] == 36497 && 
b[36498] == 36498 && 
b[36499] == 36499 && 
b[36500] == 36500 && 
b[36501] == 36501 && 
b[36502] == 36502 && 
b[36503] == 36503 && 
b[36504] == 36504 && 
b[36505] == 36505 && 
b[36506] == 36506 && 
b[36507] == 36507 && 
b[36508] == 36508 && 
b[36509] == 36509 && 
b[36510] == 36510 && 
b[36511] == 36511 && 
b[36512] == 36512 && 
b[36513] == 36513 && 
b[36514] == 36514 && 
b[36515] == 36515 && 
b[36516] == 36516 && 
b[36517] == 36517 && 
b[36518] == 36518 && 
b[36519] == 36519 && 
b[36520] == 36520 && 
b[36521] == 36521 && 
b[36522] == 36522 && 
b[36523] == 36523 && 
b[36524] == 36524 && 
b[36525] == 36525 && 
b[36526] == 36526 && 
b[36527] == 36527 && 
b[36528] == 36528 && 
b[36529] == 36529 && 
b[36530] == 36530 && 
b[36531] == 36531 && 
b[36532] == 36532 && 
b[36533] == 36533 && 
b[36534] == 36534 && 
b[36535] == 36535 && 
b[36536] == 36536 && 
b[36537] == 36537 && 
b[36538] == 36538 && 
b[36539] == 36539 && 
b[36540] == 36540 && 
b[36541] == 36541 && 
b[36542] == 36542 && 
b[36543] == 36543 && 
b[36544] == 36544 && 
b[36545] == 36545 && 
b[36546] == 36546 && 
b[36547] == 36547 && 
b[36548] == 36548 && 
b[36549] == 36549 && 
b[36550] == 36550 && 
b[36551] == 36551 && 
b[36552] == 36552 && 
b[36553] == 36553 && 
b[36554] == 36554 && 
b[36555] == 36555 && 
b[36556] == 36556 && 
b[36557] == 36557 && 
b[36558] == 36558 && 
b[36559] == 36559 && 
b[36560] == 36560 && 
b[36561] == 36561 && 
b[36562] == 36562 && 
b[36563] == 36563 && 
b[36564] == 36564 && 
b[36565] == 36565 && 
b[36566] == 36566 && 
b[36567] == 36567 && 
b[36568] == 36568 && 
b[36569] == 36569 && 
b[36570] == 36570 && 
b[36571] == 36571 && 
b[36572] == 36572 && 
b[36573] == 36573 && 
b[36574] == 36574 && 
b[36575] == 36575 && 
b[36576] == 36576 && 
b[36577] == 36577 && 
b[36578] == 36578 && 
b[36579] == 36579 && 
b[36580] == 36580 && 
b[36581] == 36581 && 
b[36582] == 36582 && 
b[36583] == 36583 && 
b[36584] == 36584 && 
b[36585] == 36585 && 
b[36586] == 36586 && 
b[36587] == 36587 && 
b[36588] == 36588 && 
b[36589] == 36589 && 
b[36590] == 36590 && 
b[36591] == 36591 && 
b[36592] == 36592 && 
b[36593] == 36593 && 
b[36594] == 36594 && 
b[36595] == 36595 && 
b[36596] == 36596 && 
b[36597] == 36597 && 
b[36598] == 36598 && 
b[36599] == 36599 && 
b[36600] == 36600 && 
b[36601] == 36601 && 
b[36602] == 36602 && 
b[36603] == 36603 && 
b[36604] == 36604 && 
b[36605] == 36605 && 
b[36606] == 36606 && 
b[36607] == 36607 && 
b[36608] == 36608 && 
b[36609] == 36609 && 
b[36610] == 36610 && 
b[36611] == 36611 && 
b[36612] == 36612 && 
b[36613] == 36613 && 
b[36614] == 36614 && 
b[36615] == 36615 && 
b[36616] == 36616 && 
b[36617] == 36617 && 
b[36618] == 36618 && 
b[36619] == 36619 && 
b[36620] == 36620 && 
b[36621] == 36621 && 
b[36622] == 36622 && 
b[36623] == 36623 && 
b[36624] == 36624 && 
b[36625] == 36625 && 
b[36626] == 36626 && 
b[36627] == 36627 && 
b[36628] == 36628 && 
b[36629] == 36629 && 
b[36630] == 36630 && 
b[36631] == 36631 && 
b[36632] == 36632 && 
b[36633] == 36633 && 
b[36634] == 36634 && 
b[36635] == 36635 && 
b[36636] == 36636 && 
b[36637] == 36637 && 
b[36638] == 36638 && 
b[36639] == 36639 && 
b[36640] == 36640 && 
b[36641] == 36641 && 
b[36642] == 36642 && 
b[36643] == 36643 && 
b[36644] == 36644 && 
b[36645] == 36645 && 
b[36646] == 36646 && 
b[36647] == 36647 && 
b[36648] == 36648 && 
b[36649] == 36649 && 
b[36650] == 36650 && 
b[36651] == 36651 && 
b[36652] == 36652 && 
b[36653] == 36653 && 
b[36654] == 36654 && 
b[36655] == 36655 && 
b[36656] == 36656 && 
b[36657] == 36657 && 
b[36658] == 36658 && 
b[36659] == 36659 && 
b[36660] == 36660 && 
b[36661] == 36661 && 
b[36662] == 36662 && 
b[36663] == 36663 && 
b[36664] == 36664 && 
b[36665] == 36665 && 
b[36666] == 36666 && 
b[36667] == 36667 && 
b[36668] == 36668 && 
b[36669] == 36669 && 
b[36670] == 36670 && 
b[36671] == 36671 && 
b[36672] == 36672 && 
b[36673] == 36673 && 
b[36674] == 36674 && 
b[36675] == 36675 && 
b[36676] == 36676 && 
b[36677] == 36677 && 
b[36678] == 36678 && 
b[36679] == 36679 && 
b[36680] == 36680 && 
b[36681] == 36681 && 
b[36682] == 36682 && 
b[36683] == 36683 && 
b[36684] == 36684 && 
b[36685] == 36685 && 
b[36686] == 36686 && 
b[36687] == 36687 && 
b[36688] == 36688 && 
b[36689] == 36689 && 
b[36690] == 36690 && 
b[36691] == 36691 && 
b[36692] == 36692 && 
b[36693] == 36693 && 
b[36694] == 36694 && 
b[36695] == 36695 && 
b[36696] == 36696 && 
b[36697] == 36697 && 
b[36698] == 36698 && 
b[36699] == 36699 && 
b[36700] == 36700 && 
b[36701] == 36701 && 
b[36702] == 36702 && 
b[36703] == 36703 && 
b[36704] == 36704 && 
b[36705] == 36705 && 
b[36706] == 36706 && 
b[36707] == 36707 && 
b[36708] == 36708 && 
b[36709] == 36709 && 
b[36710] == 36710 && 
b[36711] == 36711 && 
b[36712] == 36712 && 
b[36713] == 36713 && 
b[36714] == 36714 && 
b[36715] == 36715 && 
b[36716] == 36716 && 
b[36717] == 36717 && 
b[36718] == 36718 && 
b[36719] == 36719 && 
b[36720] == 36720 && 
b[36721] == 36721 && 
b[36722] == 36722 && 
b[36723] == 36723 && 
b[36724] == 36724 && 
b[36725] == 36725 && 
b[36726] == 36726 && 
b[36727] == 36727 && 
b[36728] == 36728 && 
b[36729] == 36729 && 
b[36730] == 36730 && 
b[36731] == 36731 && 
b[36732] == 36732 && 
b[36733] == 36733 && 
b[36734] == 36734 && 
b[36735] == 36735 && 
b[36736] == 36736 && 
b[36737] == 36737 && 
b[36738] == 36738 && 
b[36739] == 36739 && 
b[36740] == 36740 && 
b[36741] == 36741 && 
b[36742] == 36742 && 
b[36743] == 36743 && 
b[36744] == 36744 && 
b[36745] == 36745 && 
b[36746] == 36746 && 
b[36747] == 36747 && 
b[36748] == 36748 && 
b[36749] == 36749 && 
b[36750] == 36750 && 
b[36751] == 36751 && 
b[36752] == 36752 && 
b[36753] == 36753 && 
b[36754] == 36754 && 
b[36755] == 36755 && 
b[36756] == 36756 && 
b[36757] == 36757 && 
b[36758] == 36758 && 
b[36759] == 36759 && 
b[36760] == 36760 && 
b[36761] == 36761 && 
b[36762] == 36762 && 
b[36763] == 36763 && 
b[36764] == 36764 && 
b[36765] == 36765 && 
b[36766] == 36766 && 
b[36767] == 36767 && 
b[36768] == 36768 && 
b[36769] == 36769 && 
b[36770] == 36770 && 
b[36771] == 36771 && 
b[36772] == 36772 && 
b[36773] == 36773 && 
b[36774] == 36774 && 
b[36775] == 36775 && 
b[36776] == 36776 && 
b[36777] == 36777 && 
b[36778] == 36778 && 
b[36779] == 36779 && 
b[36780] == 36780 && 
b[36781] == 36781 && 
b[36782] == 36782 && 
b[36783] == 36783 && 
b[36784] == 36784 && 
b[36785] == 36785 && 
b[36786] == 36786 && 
b[36787] == 36787 && 
b[36788] == 36788 && 
b[36789] == 36789 && 
b[36790] == 36790 && 
b[36791] == 36791 && 
b[36792] == 36792 && 
b[36793] == 36793 && 
b[36794] == 36794 && 
b[36795] == 36795 && 
b[36796] == 36796 && 
b[36797] == 36797 && 
b[36798] == 36798 && 
b[36799] == 36799 && 
b[36800] == 36800 && 
b[36801] == 36801 && 
b[36802] == 36802 && 
b[36803] == 36803 && 
b[36804] == 36804 && 
b[36805] == 36805 && 
b[36806] == 36806 && 
b[36807] == 36807 && 
b[36808] == 36808 && 
b[36809] == 36809 && 
b[36810] == 36810 && 
b[36811] == 36811 && 
b[36812] == 36812 && 
b[36813] == 36813 && 
b[36814] == 36814 && 
b[36815] == 36815 && 
b[36816] == 36816 && 
b[36817] == 36817 && 
b[36818] == 36818 && 
b[36819] == 36819 && 
b[36820] == 36820 && 
b[36821] == 36821 && 
b[36822] == 36822 && 
b[36823] == 36823 && 
b[36824] == 36824 && 
b[36825] == 36825 && 
b[36826] == 36826 && 
b[36827] == 36827 && 
b[36828] == 36828 && 
b[36829] == 36829 && 
b[36830] == 36830 && 
b[36831] == 36831 && 
b[36832] == 36832 && 
b[36833] == 36833 && 
b[36834] == 36834 && 
b[36835] == 36835 && 
b[36836] == 36836 && 
b[36837] == 36837 && 
b[36838] == 36838 && 
b[36839] == 36839 && 
b[36840] == 36840 && 
b[36841] == 36841 && 
b[36842] == 36842 && 
b[36843] == 36843 && 
b[36844] == 36844 && 
b[36845] == 36845 && 
b[36846] == 36846 && 
b[36847] == 36847 && 
b[36848] == 36848 && 
b[36849] == 36849 && 
b[36850] == 36850 && 
b[36851] == 36851 && 
b[36852] == 36852 && 
b[36853] == 36853 && 
b[36854] == 36854 && 
b[36855] == 36855 && 
b[36856] == 36856 && 
b[36857] == 36857 && 
b[36858] == 36858 && 
b[36859] == 36859 && 
b[36860] == 36860 && 
b[36861] == 36861 && 
b[36862] == 36862 && 
b[36863] == 36863 && 
b[36864] == 36864 && 
b[36865] == 36865 && 
b[36866] == 36866 && 
b[36867] == 36867 && 
b[36868] == 36868 && 
b[36869] == 36869 && 
b[36870] == 36870 && 
b[36871] == 36871 && 
b[36872] == 36872 && 
b[36873] == 36873 && 
b[36874] == 36874 && 
b[36875] == 36875 && 
b[36876] == 36876 && 
b[36877] == 36877 && 
b[36878] == 36878 && 
b[36879] == 36879 && 
b[36880] == 36880 && 
b[36881] == 36881 && 
b[36882] == 36882 && 
b[36883] == 36883 && 
b[36884] == 36884 && 
b[36885] == 36885 && 
b[36886] == 36886 && 
b[36887] == 36887 && 
b[36888] == 36888 && 
b[36889] == 36889 && 
b[36890] == 36890 && 
b[36891] == 36891 && 
b[36892] == 36892 && 
b[36893] == 36893 && 
b[36894] == 36894 && 
b[36895] == 36895 && 
b[36896] == 36896 && 
b[36897] == 36897 && 
b[36898] == 36898 && 
b[36899] == 36899 && 
b[36900] == 36900 && 
b[36901] == 36901 && 
b[36902] == 36902 && 
b[36903] == 36903 && 
b[36904] == 36904 && 
b[36905] == 36905 && 
b[36906] == 36906 && 
b[36907] == 36907 && 
b[36908] == 36908 && 
b[36909] == 36909 && 
b[36910] == 36910 && 
b[36911] == 36911 && 
b[36912] == 36912 && 
b[36913] == 36913 && 
b[36914] == 36914 && 
b[36915] == 36915 && 
b[36916] == 36916 && 
b[36917] == 36917 && 
b[36918] == 36918 && 
b[36919] == 36919 && 
b[36920] == 36920 && 
b[36921] == 36921 && 
b[36922] == 36922 && 
b[36923] == 36923 && 
b[36924] == 36924 && 
b[36925] == 36925 && 
b[36926] == 36926 && 
b[36927] == 36927 && 
b[36928] == 36928 && 
b[36929] == 36929 && 
b[36930] == 36930 && 
b[36931] == 36931 && 
b[36932] == 36932 && 
b[36933] == 36933 && 
b[36934] == 36934 && 
b[36935] == 36935 && 
b[36936] == 36936 && 
b[36937] == 36937 && 
b[36938] == 36938 && 
b[36939] == 36939 && 
b[36940] == 36940 && 
b[36941] == 36941 && 
b[36942] == 36942 && 
b[36943] == 36943 && 
b[36944] == 36944 && 
b[36945] == 36945 && 
b[36946] == 36946 && 
b[36947] == 36947 && 
b[36948] == 36948 && 
b[36949] == 36949 && 
b[36950] == 36950 && 
b[36951] == 36951 && 
b[36952] == 36952 && 
b[36953] == 36953 && 
b[36954] == 36954 && 
b[36955] == 36955 && 
b[36956] == 36956 && 
b[36957] == 36957 && 
b[36958] == 36958 && 
b[36959] == 36959 && 
b[36960] == 36960 && 
b[36961] == 36961 && 
b[36962] == 36962 && 
b[36963] == 36963 && 
b[36964] == 36964 && 
b[36965] == 36965 && 
b[36966] == 36966 && 
b[36967] == 36967 && 
b[36968] == 36968 && 
b[36969] == 36969 && 
b[36970] == 36970 && 
b[36971] == 36971 && 
b[36972] == 36972 && 
b[36973] == 36973 && 
b[36974] == 36974 && 
b[36975] == 36975 && 
b[36976] == 36976 && 
b[36977] == 36977 && 
b[36978] == 36978 && 
b[36979] == 36979 && 
b[36980] == 36980 && 
b[36981] == 36981 && 
b[36982] == 36982 && 
b[36983] == 36983 && 
b[36984] == 36984 && 
b[36985] == 36985 && 
b[36986] == 36986 && 
b[36987] == 36987 && 
b[36988] == 36988 && 
b[36989] == 36989 && 
b[36990] == 36990 && 
b[36991] == 36991 && 
b[36992] == 36992 && 
b[36993] == 36993 && 
b[36994] == 36994 && 
b[36995] == 36995 && 
b[36996] == 36996 && 
b[36997] == 36997 && 
b[36998] == 36998 && 
b[36999] == 36999 && 
b[37000] == 37000 && 
b[37001] == 37001 && 
b[37002] == 37002 && 
b[37003] == 37003 && 
b[37004] == 37004 && 
b[37005] == 37005 && 
b[37006] == 37006 && 
b[37007] == 37007 && 
b[37008] == 37008 && 
b[37009] == 37009 && 
b[37010] == 37010 && 
b[37011] == 37011 && 
b[37012] == 37012 && 
b[37013] == 37013 && 
b[37014] == 37014 && 
b[37015] == 37015 && 
b[37016] == 37016 && 
b[37017] == 37017 && 
b[37018] == 37018 && 
b[37019] == 37019 && 
b[37020] == 37020 && 
b[37021] == 37021 && 
b[37022] == 37022 && 
b[37023] == 37023 && 
b[37024] == 37024 && 
b[37025] == 37025 && 
b[37026] == 37026 && 
b[37027] == 37027 && 
b[37028] == 37028 && 
b[37029] == 37029 && 
b[37030] == 37030 && 
b[37031] == 37031 && 
b[37032] == 37032 && 
b[37033] == 37033 && 
b[37034] == 37034 && 
b[37035] == 37035 && 
b[37036] == 37036 && 
b[37037] == 37037 && 
b[37038] == 37038 && 
b[37039] == 37039 && 
b[37040] == 37040 && 
b[37041] == 37041 && 
b[37042] == 37042 && 
b[37043] == 37043 && 
b[37044] == 37044 && 
b[37045] == 37045 && 
b[37046] == 37046 && 
b[37047] == 37047 && 
b[37048] == 37048 && 
b[37049] == 37049 && 
b[37050] == 37050 && 
b[37051] == 37051 && 
b[37052] == 37052 && 
b[37053] == 37053 && 
b[37054] == 37054 && 
b[37055] == 37055 && 
b[37056] == 37056 && 
b[37057] == 37057 && 
b[37058] == 37058 && 
b[37059] == 37059 && 
b[37060] == 37060 && 
b[37061] == 37061 && 
b[37062] == 37062 && 
b[37063] == 37063 && 
b[37064] == 37064 && 
b[37065] == 37065 && 
b[37066] == 37066 && 
b[37067] == 37067 && 
b[37068] == 37068 && 
b[37069] == 37069 && 
b[37070] == 37070 && 
b[37071] == 37071 && 
b[37072] == 37072 && 
b[37073] == 37073 && 
b[37074] == 37074 && 
b[37075] == 37075 && 
b[37076] == 37076 && 
b[37077] == 37077 && 
b[37078] == 37078 && 
b[37079] == 37079 && 
b[37080] == 37080 && 
b[37081] == 37081 && 
b[37082] == 37082 && 
b[37083] == 37083 && 
b[37084] == 37084 && 
b[37085] == 37085 && 
b[37086] == 37086 && 
b[37087] == 37087 && 
b[37088] == 37088 && 
b[37089] == 37089 && 
b[37090] == 37090 && 
b[37091] == 37091 && 
b[37092] == 37092 && 
b[37093] == 37093 && 
b[37094] == 37094 && 
b[37095] == 37095 && 
b[37096] == 37096 && 
b[37097] == 37097 && 
b[37098] == 37098 && 
b[37099] == 37099 && 
b[37100] == 37100 && 
b[37101] == 37101 && 
b[37102] == 37102 && 
b[37103] == 37103 && 
b[37104] == 37104 && 
b[37105] == 37105 && 
b[37106] == 37106 && 
b[37107] == 37107 && 
b[37108] == 37108 && 
b[37109] == 37109 && 
b[37110] == 37110 && 
b[37111] == 37111 && 
b[37112] == 37112 && 
b[37113] == 37113 && 
b[37114] == 37114 && 
b[37115] == 37115 && 
b[37116] == 37116 && 
b[37117] == 37117 && 
b[37118] == 37118 && 
b[37119] == 37119 && 
b[37120] == 37120 && 
b[37121] == 37121 && 
b[37122] == 37122 && 
b[37123] == 37123 && 
b[37124] == 37124 && 
b[37125] == 37125 && 
b[37126] == 37126 && 
b[37127] == 37127 && 
b[37128] == 37128 && 
b[37129] == 37129 && 
b[37130] == 37130 && 
b[37131] == 37131 && 
b[37132] == 37132 && 
b[37133] == 37133 && 
b[37134] == 37134 && 
b[37135] == 37135 && 
b[37136] == 37136 && 
b[37137] == 37137 && 
b[37138] == 37138 && 
b[37139] == 37139 && 
b[37140] == 37140 && 
b[37141] == 37141 && 
b[37142] == 37142 && 
b[37143] == 37143 && 
b[37144] == 37144 && 
b[37145] == 37145 && 
b[37146] == 37146 && 
b[37147] == 37147 && 
b[37148] == 37148 && 
b[37149] == 37149 && 
b[37150] == 37150 && 
b[37151] == 37151 && 
b[37152] == 37152 && 
b[37153] == 37153 && 
b[37154] == 37154 && 
b[37155] == 37155 && 
b[37156] == 37156 && 
b[37157] == 37157 && 
b[37158] == 37158 && 
b[37159] == 37159 && 
b[37160] == 37160 && 
b[37161] == 37161 && 
b[37162] == 37162 && 
b[37163] == 37163 && 
b[37164] == 37164 && 
b[37165] == 37165 && 
b[37166] == 37166 && 
b[37167] == 37167 && 
b[37168] == 37168 && 
b[37169] == 37169 && 
b[37170] == 37170 && 
b[37171] == 37171 && 
b[37172] == 37172 && 
b[37173] == 37173 && 
b[37174] == 37174 && 
b[37175] == 37175 && 
b[37176] == 37176 && 
b[37177] == 37177 && 
b[37178] == 37178 && 
b[37179] == 37179 && 
b[37180] == 37180 && 
b[37181] == 37181 && 
b[37182] == 37182 && 
b[37183] == 37183 && 
b[37184] == 37184 && 
b[37185] == 37185 && 
b[37186] == 37186 && 
b[37187] == 37187 && 
b[37188] == 37188 && 
b[37189] == 37189 && 
b[37190] == 37190 && 
b[37191] == 37191 && 
b[37192] == 37192 && 
b[37193] == 37193 && 
b[37194] == 37194 && 
b[37195] == 37195 && 
b[37196] == 37196 && 
b[37197] == 37197 && 
b[37198] == 37198 && 
b[37199] == 37199 && 
b[37200] == 37200 && 
b[37201] == 37201 && 
b[37202] == 37202 && 
b[37203] == 37203 && 
b[37204] == 37204 && 
b[37205] == 37205 && 
b[37206] == 37206 && 
b[37207] == 37207 && 
b[37208] == 37208 && 
b[37209] == 37209 && 
b[37210] == 37210 && 
b[37211] == 37211 && 
b[37212] == 37212 && 
b[37213] == 37213 && 
b[37214] == 37214 && 
b[37215] == 37215 && 
b[37216] == 37216 && 
b[37217] == 37217 && 
b[37218] == 37218 && 
b[37219] == 37219 && 
b[37220] == 37220 && 
b[37221] == 37221 && 
b[37222] == 37222 && 
b[37223] == 37223 && 
b[37224] == 37224 && 
b[37225] == 37225 && 
b[37226] == 37226 && 
b[37227] == 37227 && 
b[37228] == 37228 && 
b[37229] == 37229 && 
b[37230] == 37230 && 
b[37231] == 37231 && 
b[37232] == 37232 && 
b[37233] == 37233 && 
b[37234] == 37234 && 
b[37235] == 37235 && 
b[37236] == 37236 && 
b[37237] == 37237 && 
b[37238] == 37238 && 
b[37239] == 37239 && 
b[37240] == 37240 && 
b[37241] == 37241 && 
b[37242] == 37242 && 
b[37243] == 37243 && 
b[37244] == 37244 && 
b[37245] == 37245 && 
b[37246] == 37246 && 
b[37247] == 37247 && 
b[37248] == 37248 && 
b[37249] == 37249 && 
b[37250] == 37250 && 
b[37251] == 37251 && 
b[37252] == 37252 && 
b[37253] == 37253 && 
b[37254] == 37254 && 
b[37255] == 37255 && 
b[37256] == 37256 && 
b[37257] == 37257 && 
b[37258] == 37258 && 
b[37259] == 37259 && 
b[37260] == 37260 && 
b[37261] == 37261 && 
b[37262] == 37262 && 
b[37263] == 37263 && 
b[37264] == 37264 && 
b[37265] == 37265 && 
b[37266] == 37266 && 
b[37267] == 37267 && 
b[37268] == 37268 && 
b[37269] == 37269 && 
b[37270] == 37270 && 
b[37271] == 37271 && 
b[37272] == 37272 && 
b[37273] == 37273 && 
b[37274] == 37274 && 
b[37275] == 37275 && 
b[37276] == 37276 && 
b[37277] == 37277 && 
b[37278] == 37278 && 
b[37279] == 37279 && 
b[37280] == 37280 && 
b[37281] == 37281 && 
b[37282] == 37282 && 
b[37283] == 37283 && 
b[37284] == 37284 && 
b[37285] == 37285 && 
b[37286] == 37286 && 
b[37287] == 37287 && 
b[37288] == 37288 && 
b[37289] == 37289 && 
b[37290] == 37290 && 
b[37291] == 37291 && 
b[37292] == 37292 && 
b[37293] == 37293 && 
b[37294] == 37294 && 
b[37295] == 37295 && 
b[37296] == 37296 && 
b[37297] == 37297 && 
b[37298] == 37298 && 
b[37299] == 37299 && 
b[37300] == 37300 && 
b[37301] == 37301 && 
b[37302] == 37302 && 
b[37303] == 37303 && 
b[37304] == 37304 && 
b[37305] == 37305 && 
b[37306] == 37306 && 
b[37307] == 37307 && 
b[37308] == 37308 && 
b[37309] == 37309 && 
b[37310] == 37310 && 
b[37311] == 37311 && 
b[37312] == 37312 && 
b[37313] == 37313 && 
b[37314] == 37314 && 
b[37315] == 37315 && 
b[37316] == 37316 && 
b[37317] == 37317 && 
b[37318] == 37318 && 
b[37319] == 37319 && 
b[37320] == 37320 && 
b[37321] == 37321 && 
b[37322] == 37322 && 
b[37323] == 37323 && 
b[37324] == 37324 && 
b[37325] == 37325 && 
b[37326] == 37326 && 
b[37327] == 37327 && 
b[37328] == 37328 && 
b[37329] == 37329 && 
b[37330] == 37330 && 
b[37331] == 37331 && 
b[37332] == 37332 && 
b[37333] == 37333 && 
b[37334] == 37334 && 
b[37335] == 37335 && 
b[37336] == 37336 && 
b[37337] == 37337 && 
b[37338] == 37338 && 
b[37339] == 37339 && 
b[37340] == 37340 && 
b[37341] == 37341 && 
b[37342] == 37342 && 
b[37343] == 37343 && 
b[37344] == 37344 && 
b[37345] == 37345 && 
b[37346] == 37346 && 
b[37347] == 37347 && 
b[37348] == 37348 && 
b[37349] == 37349 && 
b[37350] == 37350 && 
b[37351] == 37351 && 
b[37352] == 37352 && 
b[37353] == 37353 && 
b[37354] == 37354 && 
b[37355] == 37355 && 
b[37356] == 37356 && 
b[37357] == 37357 && 
b[37358] == 37358 && 
b[37359] == 37359 && 
b[37360] == 37360 && 
b[37361] == 37361 && 
b[37362] == 37362 && 
b[37363] == 37363 && 
b[37364] == 37364 && 
b[37365] == 37365 && 
b[37366] == 37366 && 
b[37367] == 37367 && 
b[37368] == 37368 && 
b[37369] == 37369 && 
b[37370] == 37370 && 
b[37371] == 37371 && 
b[37372] == 37372 && 
b[37373] == 37373 && 
b[37374] == 37374 && 
b[37375] == 37375 && 
b[37376] == 37376 && 
b[37377] == 37377 && 
b[37378] == 37378 && 
b[37379] == 37379 && 
b[37380] == 37380 && 
b[37381] == 37381 && 
b[37382] == 37382 && 
b[37383] == 37383 && 
b[37384] == 37384 && 
b[37385] == 37385 && 
b[37386] == 37386 && 
b[37387] == 37387 && 
b[37388] == 37388 && 
b[37389] == 37389 && 
b[37390] == 37390 && 
b[37391] == 37391 && 
b[37392] == 37392 && 
b[37393] == 37393 && 
b[37394] == 37394 && 
b[37395] == 37395 && 
b[37396] == 37396 && 
b[37397] == 37397 && 
b[37398] == 37398 && 
b[37399] == 37399 && 
b[37400] == 37400 && 
b[37401] == 37401 && 
b[37402] == 37402 && 
b[37403] == 37403 && 
b[37404] == 37404 && 
b[37405] == 37405 && 
b[37406] == 37406 && 
b[37407] == 37407 && 
b[37408] == 37408 && 
b[37409] == 37409 && 
b[37410] == 37410 && 
b[37411] == 37411 && 
b[37412] == 37412 && 
b[37413] == 37413 && 
b[37414] == 37414 && 
b[37415] == 37415 && 
b[37416] == 37416 && 
b[37417] == 37417 && 
b[37418] == 37418 && 
b[37419] == 37419 && 
b[37420] == 37420 && 
b[37421] == 37421 && 
b[37422] == 37422 && 
b[37423] == 37423 && 
b[37424] == 37424 && 
b[37425] == 37425 && 
b[37426] == 37426 && 
b[37427] == 37427 && 
b[37428] == 37428 && 
b[37429] == 37429 && 
b[37430] == 37430 && 
b[37431] == 37431 && 
b[37432] == 37432 && 
b[37433] == 37433 && 
b[37434] == 37434 && 
b[37435] == 37435 && 
b[37436] == 37436 && 
b[37437] == 37437 && 
b[37438] == 37438 && 
b[37439] == 37439 && 
b[37440] == 37440 && 
b[37441] == 37441 && 
b[37442] == 37442 && 
b[37443] == 37443 && 
b[37444] == 37444 && 
b[37445] == 37445 && 
b[37446] == 37446 && 
b[37447] == 37447 && 
b[37448] == 37448 && 
b[37449] == 37449 && 
b[37450] == 37450 && 
b[37451] == 37451 && 
b[37452] == 37452 && 
b[37453] == 37453 && 
b[37454] == 37454 && 
b[37455] == 37455 && 
b[37456] == 37456 && 
b[37457] == 37457 && 
b[37458] == 37458 && 
b[37459] == 37459 && 
b[37460] == 37460 && 
b[37461] == 37461 && 
b[37462] == 37462 && 
b[37463] == 37463 && 
b[37464] == 37464 && 
b[37465] == 37465 && 
b[37466] == 37466 && 
b[37467] == 37467 && 
b[37468] == 37468 && 
b[37469] == 37469 && 
b[37470] == 37470 && 
b[37471] == 37471 && 
b[37472] == 37472 && 
b[37473] == 37473 && 
b[37474] == 37474 && 
b[37475] == 37475 && 
b[37476] == 37476 && 
b[37477] == 37477 && 
b[37478] == 37478 && 
b[37479] == 37479 && 
b[37480] == 37480 && 
b[37481] == 37481 && 
b[37482] == 37482 && 
b[37483] == 37483 && 
b[37484] == 37484 && 
b[37485] == 37485 && 
b[37486] == 37486 && 
b[37487] == 37487 && 
b[37488] == 37488 && 
b[37489] == 37489 && 
b[37490] == 37490 && 
b[37491] == 37491 && 
b[37492] == 37492 && 
b[37493] == 37493 && 
b[37494] == 37494 && 
b[37495] == 37495 && 
b[37496] == 37496 && 
b[37497] == 37497 && 
b[37498] == 37498 && 
b[37499] == 37499 && 
b[37500] == 37500 && 
b[37501] == 37501 && 
b[37502] == 37502 && 
b[37503] == 37503 && 
b[37504] == 37504 && 
b[37505] == 37505 && 
b[37506] == 37506 && 
b[37507] == 37507 && 
b[37508] == 37508 && 
b[37509] == 37509 && 
b[37510] == 37510 && 
b[37511] == 37511 && 
b[37512] == 37512 && 
b[37513] == 37513 && 
b[37514] == 37514 && 
b[37515] == 37515 && 
b[37516] == 37516 && 
b[37517] == 37517 && 
b[37518] == 37518 && 
b[37519] == 37519 && 
b[37520] == 37520 && 
b[37521] == 37521 && 
b[37522] == 37522 && 
b[37523] == 37523 && 
b[37524] == 37524 && 
b[37525] == 37525 && 
b[37526] == 37526 && 
b[37527] == 37527 && 
b[37528] == 37528 && 
b[37529] == 37529 && 
b[37530] == 37530 && 
b[37531] == 37531 && 
b[37532] == 37532 && 
b[37533] == 37533 && 
b[37534] == 37534 && 
b[37535] == 37535 && 
b[37536] == 37536 && 
b[37537] == 37537 && 
b[37538] == 37538 && 
b[37539] == 37539 && 
b[37540] == 37540 && 
b[37541] == 37541 && 
b[37542] == 37542 && 
b[37543] == 37543 && 
b[37544] == 37544 && 
b[37545] == 37545 && 
b[37546] == 37546 && 
b[37547] == 37547 && 
b[37548] == 37548 && 
b[37549] == 37549 && 
b[37550] == 37550 && 
b[37551] == 37551 && 
b[37552] == 37552 && 
b[37553] == 37553 && 
b[37554] == 37554 && 
b[37555] == 37555 && 
b[37556] == 37556 && 
b[37557] == 37557 && 
b[37558] == 37558 && 
b[37559] == 37559 && 
b[37560] == 37560 && 
b[37561] == 37561 && 
b[37562] == 37562 && 
b[37563] == 37563 && 
b[37564] == 37564 && 
b[37565] == 37565 && 
b[37566] == 37566 && 
b[37567] == 37567 && 
b[37568] == 37568 && 
b[37569] == 37569 && 
b[37570] == 37570 && 
b[37571] == 37571 && 
b[37572] == 37572 && 
b[37573] == 37573 && 
b[37574] == 37574 && 
b[37575] == 37575 && 
b[37576] == 37576 && 
b[37577] == 37577 && 
b[37578] == 37578 && 
b[37579] == 37579 && 
b[37580] == 37580 && 
b[37581] == 37581 && 
b[37582] == 37582 && 
b[37583] == 37583 && 
b[37584] == 37584 && 
b[37585] == 37585 && 
b[37586] == 37586 && 
b[37587] == 37587 && 
b[37588] == 37588 && 
b[37589] == 37589 && 
b[37590] == 37590 && 
b[37591] == 37591 && 
b[37592] == 37592 && 
b[37593] == 37593 && 
b[37594] == 37594 && 
b[37595] == 37595 && 
b[37596] == 37596 && 
b[37597] == 37597 && 
b[37598] == 37598 && 
b[37599] == 37599 && 
b[37600] == 37600 && 
b[37601] == 37601 && 
b[37602] == 37602 && 
b[37603] == 37603 && 
b[37604] == 37604 && 
b[37605] == 37605 && 
b[37606] == 37606 && 
b[37607] == 37607 && 
b[37608] == 37608 && 
b[37609] == 37609 && 
b[37610] == 37610 && 
b[37611] == 37611 && 
b[37612] == 37612 && 
b[37613] == 37613 && 
b[37614] == 37614 && 
b[37615] == 37615 && 
b[37616] == 37616 && 
b[37617] == 37617 && 
b[37618] == 37618 && 
b[37619] == 37619 && 
b[37620] == 37620 && 
b[37621] == 37621 && 
b[37622] == 37622 && 
b[37623] == 37623 && 
b[37624] == 37624 && 
b[37625] == 37625 && 
b[37626] == 37626 && 
b[37627] == 37627 && 
b[37628] == 37628 && 
b[37629] == 37629 && 
b[37630] == 37630 && 
b[37631] == 37631 && 
b[37632] == 37632 && 
b[37633] == 37633 && 
b[37634] == 37634 && 
b[37635] == 37635 && 
b[37636] == 37636 && 
b[37637] == 37637 && 
b[37638] == 37638 && 
b[37639] == 37639 && 
b[37640] == 37640 && 
b[37641] == 37641 && 
b[37642] == 37642 && 
b[37643] == 37643 && 
b[37644] == 37644 && 
b[37645] == 37645 && 
b[37646] == 37646 && 
b[37647] == 37647 && 
b[37648] == 37648 && 
b[37649] == 37649 && 
b[37650] == 37650 && 
b[37651] == 37651 && 
b[37652] == 37652 && 
b[37653] == 37653 && 
b[37654] == 37654 && 
b[37655] == 37655 && 
b[37656] == 37656 && 
b[37657] == 37657 && 
b[37658] == 37658 && 
b[37659] == 37659 && 
b[37660] == 37660 && 
b[37661] == 37661 && 
b[37662] == 37662 && 
b[37663] == 37663 && 
b[37664] == 37664 && 
b[37665] == 37665 && 
b[37666] == 37666 && 
b[37667] == 37667 && 
b[37668] == 37668 && 
b[37669] == 37669 && 
b[37670] == 37670 && 
b[37671] == 37671 && 
b[37672] == 37672 && 
b[37673] == 37673 && 
b[37674] == 37674 && 
b[37675] == 37675 && 
b[37676] == 37676 && 
b[37677] == 37677 && 
b[37678] == 37678 && 
b[37679] == 37679 && 
b[37680] == 37680 && 
b[37681] == 37681 && 
b[37682] == 37682 && 
b[37683] == 37683 && 
b[37684] == 37684 && 
b[37685] == 37685 && 
b[37686] == 37686 && 
b[37687] == 37687 && 
b[37688] == 37688 && 
b[37689] == 37689 && 
b[37690] == 37690 && 
b[37691] == 37691 && 
b[37692] == 37692 && 
b[37693] == 37693 && 
b[37694] == 37694 && 
b[37695] == 37695 && 
b[37696] == 37696 && 
b[37697] == 37697 && 
b[37698] == 37698 && 
b[37699] == 37699 && 
b[37700] == 37700 && 
b[37701] == 37701 && 
b[37702] == 37702 && 
b[37703] == 37703 && 
b[37704] == 37704 && 
b[37705] == 37705 && 
b[37706] == 37706 && 
b[37707] == 37707 && 
b[37708] == 37708 && 
b[37709] == 37709 && 
b[37710] == 37710 && 
b[37711] == 37711 && 
b[37712] == 37712 && 
b[37713] == 37713 && 
b[37714] == 37714 && 
b[37715] == 37715 && 
b[37716] == 37716 && 
b[37717] == 37717 && 
b[37718] == 37718 && 
b[37719] == 37719 && 
b[37720] == 37720 && 
b[37721] == 37721 && 
b[37722] == 37722 && 
b[37723] == 37723 && 
b[37724] == 37724 && 
b[37725] == 37725 && 
b[37726] == 37726 && 
b[37727] == 37727 && 
b[37728] == 37728 && 
b[37729] == 37729 && 
b[37730] == 37730 && 
b[37731] == 37731 && 
b[37732] == 37732 && 
b[37733] == 37733 && 
b[37734] == 37734 && 
b[37735] == 37735 && 
b[37736] == 37736 && 
b[37737] == 37737 && 
b[37738] == 37738 && 
b[37739] == 37739 && 
b[37740] == 37740 && 
b[37741] == 37741 && 
b[37742] == 37742 && 
b[37743] == 37743 && 
b[37744] == 37744 && 
b[37745] == 37745 && 
b[37746] == 37746 && 
b[37747] == 37747 && 
b[37748] == 37748 && 
b[37749] == 37749 && 
b[37750] == 37750 && 
b[37751] == 37751 && 
b[37752] == 37752 && 
b[37753] == 37753 && 
b[37754] == 37754 && 
b[37755] == 37755 && 
b[37756] == 37756 && 
b[37757] == 37757 && 
b[37758] == 37758 && 
b[37759] == 37759 && 
b[37760] == 37760 && 
b[37761] == 37761 && 
b[37762] == 37762 && 
b[37763] == 37763 && 
b[37764] == 37764 && 
b[37765] == 37765 && 
b[37766] == 37766 && 
b[37767] == 37767 && 
b[37768] == 37768 && 
b[37769] == 37769 && 
b[37770] == 37770 && 
b[37771] == 37771 && 
b[37772] == 37772 && 
b[37773] == 37773 && 
b[37774] == 37774 && 
b[37775] == 37775 && 
b[37776] == 37776 && 
b[37777] == 37777 && 
b[37778] == 37778 && 
b[37779] == 37779 && 
b[37780] == 37780 && 
b[37781] == 37781 && 
b[37782] == 37782 && 
b[37783] == 37783 && 
b[37784] == 37784 && 
b[37785] == 37785 && 
b[37786] == 37786 && 
b[37787] == 37787 && 
b[37788] == 37788 && 
b[37789] == 37789 && 
b[37790] == 37790 && 
b[37791] == 37791 && 
b[37792] == 37792 && 
b[37793] == 37793 && 
b[37794] == 37794 && 
b[37795] == 37795 && 
b[37796] == 37796 && 
b[37797] == 37797 && 
b[37798] == 37798 && 
b[37799] == 37799 && 
b[37800] == 37800 && 
b[37801] == 37801 && 
b[37802] == 37802 && 
b[37803] == 37803 && 
b[37804] == 37804 && 
b[37805] == 37805 && 
b[37806] == 37806 && 
b[37807] == 37807 && 
b[37808] == 37808 && 
b[37809] == 37809 && 
b[37810] == 37810 && 
b[37811] == 37811 && 
b[37812] == 37812 && 
b[37813] == 37813 && 
b[37814] == 37814 && 
b[37815] == 37815 && 
b[37816] == 37816 && 
b[37817] == 37817 && 
b[37818] == 37818 && 
b[37819] == 37819 && 
b[37820] == 37820 && 
b[37821] == 37821 && 
b[37822] == 37822 && 
b[37823] == 37823 && 
b[37824] == 37824 && 
b[37825] == 37825 && 
b[37826] == 37826 && 
b[37827] == 37827 && 
b[37828] == 37828 && 
b[37829] == 37829 && 
b[37830] == 37830 && 
b[37831] == 37831 && 
b[37832] == 37832 && 
b[37833] == 37833 && 
b[37834] == 37834 && 
b[37835] == 37835 && 
b[37836] == 37836 && 
b[37837] == 37837 && 
b[37838] == 37838 && 
b[37839] == 37839 && 
b[37840] == 37840 && 
b[37841] == 37841 && 
b[37842] == 37842 && 
b[37843] == 37843 && 
b[37844] == 37844 && 
b[37845] == 37845 && 
b[37846] == 37846 && 
b[37847] == 37847 && 
b[37848] == 37848 && 
b[37849] == 37849 && 
b[37850] == 37850 && 
b[37851] == 37851 && 
b[37852] == 37852 && 
b[37853] == 37853 && 
b[37854] == 37854 && 
b[37855] == 37855 && 
b[37856] == 37856 && 
b[37857] == 37857 && 
b[37858] == 37858 && 
b[37859] == 37859 && 
b[37860] == 37860 && 
b[37861] == 37861 && 
b[37862] == 37862 && 
b[37863] == 37863 && 
b[37864] == 37864 && 
b[37865] == 37865 && 
b[37866] == 37866 && 
b[37867] == 37867 && 
b[37868] == 37868 && 
b[37869] == 37869 && 
b[37870] == 37870 && 
b[37871] == 37871 && 
b[37872] == 37872 && 
b[37873] == 37873 && 
b[37874] == 37874 && 
b[37875] == 37875 && 
b[37876] == 37876 && 
b[37877] == 37877 && 
b[37878] == 37878 && 
b[37879] == 37879 && 
b[37880] == 37880 && 
b[37881] == 37881 && 
b[37882] == 37882 && 
b[37883] == 37883 && 
b[37884] == 37884 && 
b[37885] == 37885 && 
b[37886] == 37886 && 
b[37887] == 37887 && 
b[37888] == 37888 && 
b[37889] == 37889 && 
b[37890] == 37890 && 
b[37891] == 37891 && 
b[37892] == 37892 && 
b[37893] == 37893 && 
b[37894] == 37894 && 
b[37895] == 37895 && 
b[37896] == 37896 && 
b[37897] == 37897 && 
b[37898] == 37898 && 
b[37899] == 37899 && 
b[37900] == 37900 && 
b[37901] == 37901 && 
b[37902] == 37902 && 
b[37903] == 37903 && 
b[37904] == 37904 && 
b[37905] == 37905 && 
b[37906] == 37906 && 
b[37907] == 37907 && 
b[37908] == 37908 && 
b[37909] == 37909 && 
b[37910] == 37910 && 
b[37911] == 37911 && 
b[37912] == 37912 && 
b[37913] == 37913 && 
b[37914] == 37914 && 
b[37915] == 37915 && 
b[37916] == 37916 && 
b[37917] == 37917 && 
b[37918] == 37918 && 
b[37919] == 37919 && 
b[37920] == 37920 && 
b[37921] == 37921 && 
b[37922] == 37922 && 
b[37923] == 37923 && 
b[37924] == 37924 && 
b[37925] == 37925 && 
b[37926] == 37926 && 
b[37927] == 37927 && 
b[37928] == 37928 && 
b[37929] == 37929 && 
b[37930] == 37930 && 
b[37931] == 37931 && 
b[37932] == 37932 && 
b[37933] == 37933 && 
b[37934] == 37934 && 
b[37935] == 37935 && 
b[37936] == 37936 && 
b[37937] == 37937 && 
b[37938] == 37938 && 
b[37939] == 37939 && 
b[37940] == 37940 && 
b[37941] == 37941 && 
b[37942] == 37942 && 
b[37943] == 37943 && 
b[37944] == 37944 && 
b[37945] == 37945 && 
b[37946] == 37946 && 
b[37947] == 37947 && 
b[37948] == 37948 && 
b[37949] == 37949 && 
b[37950] == 37950 && 
b[37951] == 37951 && 
b[37952] == 37952 && 
b[37953] == 37953 && 
b[37954] == 37954 && 
b[37955] == 37955 && 
b[37956] == 37956 && 
b[37957] == 37957 && 
b[37958] == 37958 && 
b[37959] == 37959 && 
b[37960] == 37960 && 
b[37961] == 37961 && 
b[37962] == 37962 && 
b[37963] == 37963 && 
b[37964] == 37964 && 
b[37965] == 37965 && 
b[37966] == 37966 && 
b[37967] == 37967 && 
b[37968] == 37968 && 
b[37969] == 37969 && 
b[37970] == 37970 && 
b[37971] == 37971 && 
b[37972] == 37972 && 
b[37973] == 37973 && 
b[37974] == 37974 && 
b[37975] == 37975 && 
b[37976] == 37976 && 
b[37977] == 37977 && 
b[37978] == 37978 && 
b[37979] == 37979 && 
b[37980] == 37980 && 
b[37981] == 37981 && 
b[37982] == 37982 && 
b[37983] == 37983 && 
b[37984] == 37984 && 
b[37985] == 37985 && 
b[37986] == 37986 && 
b[37987] == 37987 && 
b[37988] == 37988 && 
b[37989] == 37989 && 
b[37990] == 37990 && 
b[37991] == 37991 && 
b[37992] == 37992 && 
b[37993] == 37993 && 
b[37994] == 37994 && 
b[37995] == 37995 && 
b[37996] == 37996 && 
b[37997] == 37997 && 
b[37998] == 37998 && 
b[37999] == 37999 && 
b[38000] == 38000 && 
b[38001] == 38001 && 
b[38002] == 38002 && 
b[38003] == 38003 && 
b[38004] == 38004 && 
b[38005] == 38005 && 
b[38006] == 38006 && 
b[38007] == 38007 && 
b[38008] == 38008 && 
b[38009] == 38009 && 
b[38010] == 38010 && 
b[38011] == 38011 && 
b[38012] == 38012 && 
b[38013] == 38013 && 
b[38014] == 38014 && 
b[38015] == 38015 && 
b[38016] == 38016 && 
b[38017] == 38017 && 
b[38018] == 38018 && 
b[38019] == 38019 && 
b[38020] == 38020 && 
b[38021] == 38021 && 
b[38022] == 38022 && 
b[38023] == 38023 && 
b[38024] == 38024 && 
b[38025] == 38025 && 
b[38026] == 38026 && 
b[38027] == 38027 && 
b[38028] == 38028 && 
b[38029] == 38029 && 
b[38030] == 38030 && 
b[38031] == 38031 && 
b[38032] == 38032 && 
b[38033] == 38033 && 
b[38034] == 38034 && 
b[38035] == 38035 && 
b[38036] == 38036 && 
b[38037] == 38037 && 
b[38038] == 38038 && 
b[38039] == 38039 && 
b[38040] == 38040 && 
b[38041] == 38041 && 
b[38042] == 38042 && 
b[38043] == 38043 && 
b[38044] == 38044 && 
b[38045] == 38045 && 
b[38046] == 38046 && 
b[38047] == 38047 && 
b[38048] == 38048 && 
b[38049] == 38049 && 
b[38050] == 38050 && 
b[38051] == 38051 && 
b[38052] == 38052 && 
b[38053] == 38053 && 
b[38054] == 38054 && 
b[38055] == 38055 && 
b[38056] == 38056 && 
b[38057] == 38057 && 
b[38058] == 38058 && 
b[38059] == 38059 && 
b[38060] == 38060 && 
b[38061] == 38061 && 
b[38062] == 38062 && 
b[38063] == 38063 && 
b[38064] == 38064 && 
b[38065] == 38065 && 
b[38066] == 38066 && 
b[38067] == 38067 && 
b[38068] == 38068 && 
b[38069] == 38069 && 
b[38070] == 38070 && 
b[38071] == 38071 && 
b[38072] == 38072 && 
b[38073] == 38073 && 
b[38074] == 38074 && 
b[38075] == 38075 && 
b[38076] == 38076 && 
b[38077] == 38077 && 
b[38078] == 38078 && 
b[38079] == 38079 && 
b[38080] == 38080 && 
b[38081] == 38081 && 
b[38082] == 38082 && 
b[38083] == 38083 && 
b[38084] == 38084 && 
b[38085] == 38085 && 
b[38086] == 38086 && 
b[38087] == 38087 && 
b[38088] == 38088 && 
b[38089] == 38089 && 
b[38090] == 38090 && 
b[38091] == 38091 && 
b[38092] == 38092 && 
b[38093] == 38093 && 
b[38094] == 38094 && 
b[38095] == 38095 && 
b[38096] == 38096 && 
b[38097] == 38097 && 
b[38098] == 38098 && 
b[38099] == 38099 && 
b[38100] == 38100 && 
b[38101] == 38101 && 
b[38102] == 38102 && 
b[38103] == 38103 && 
b[38104] == 38104 && 
b[38105] == 38105 && 
b[38106] == 38106 && 
b[38107] == 38107 && 
b[38108] == 38108 && 
b[38109] == 38109 && 
b[38110] == 38110 && 
b[38111] == 38111 && 
b[38112] == 38112 && 
b[38113] == 38113 && 
b[38114] == 38114 && 
b[38115] == 38115 && 
b[38116] == 38116 && 
b[38117] == 38117 && 
b[38118] == 38118 && 
b[38119] == 38119 && 
b[38120] == 38120 && 
b[38121] == 38121 && 
b[38122] == 38122 && 
b[38123] == 38123 && 
b[38124] == 38124 && 
b[38125] == 38125 && 
b[38126] == 38126 && 
b[38127] == 38127 && 
b[38128] == 38128 && 
b[38129] == 38129 && 
b[38130] == 38130 && 
b[38131] == 38131 && 
b[38132] == 38132 && 
b[38133] == 38133 && 
b[38134] == 38134 && 
b[38135] == 38135 && 
b[38136] == 38136 && 
b[38137] == 38137 && 
b[38138] == 38138 && 
b[38139] == 38139 && 
b[38140] == 38140 && 
b[38141] == 38141 && 
b[38142] == 38142 && 
b[38143] == 38143 && 
b[38144] == 38144 && 
b[38145] == 38145 && 
b[38146] == 38146 && 
b[38147] == 38147 && 
b[38148] == 38148 && 
b[38149] == 38149 && 
b[38150] == 38150 && 
b[38151] == 38151 && 
b[38152] == 38152 && 
b[38153] == 38153 && 
b[38154] == 38154 && 
b[38155] == 38155 && 
b[38156] == 38156 && 
b[38157] == 38157 && 
b[38158] == 38158 && 
b[38159] == 38159 && 
b[38160] == 38160 && 
b[38161] == 38161 && 
b[38162] == 38162 && 
b[38163] == 38163 && 
b[38164] == 38164 && 
b[38165] == 38165 && 
b[38166] == 38166 && 
b[38167] == 38167 && 
b[38168] == 38168 && 
b[38169] == 38169 && 
b[38170] == 38170 && 
b[38171] == 38171 && 
b[38172] == 38172 && 
b[38173] == 38173 && 
b[38174] == 38174 && 
b[38175] == 38175 && 
b[38176] == 38176 && 
b[38177] == 38177 && 
b[38178] == 38178 && 
b[38179] == 38179 && 
b[38180] == 38180 && 
b[38181] == 38181 && 
b[38182] == 38182 && 
b[38183] == 38183 && 
b[38184] == 38184 && 
b[38185] == 38185 && 
b[38186] == 38186 && 
b[38187] == 38187 && 
b[38188] == 38188 && 
b[38189] == 38189 && 
b[38190] == 38190 && 
b[38191] == 38191 && 
b[38192] == 38192 && 
b[38193] == 38193 && 
b[38194] == 38194 && 
b[38195] == 38195 && 
b[38196] == 38196 && 
b[38197] == 38197 && 
b[38198] == 38198 && 
b[38199] == 38199 && 
b[38200] == 38200 && 
b[38201] == 38201 && 
b[38202] == 38202 && 
b[38203] == 38203 && 
b[38204] == 38204 && 
b[38205] == 38205 && 
b[38206] == 38206 && 
b[38207] == 38207 && 
b[38208] == 38208 && 
b[38209] == 38209 && 
b[38210] == 38210 && 
b[38211] == 38211 && 
b[38212] == 38212 && 
b[38213] == 38213 && 
b[38214] == 38214 && 
b[38215] == 38215 && 
b[38216] == 38216 && 
b[38217] == 38217 && 
b[38218] == 38218 && 
b[38219] == 38219 && 
b[38220] == 38220 && 
b[38221] == 38221 && 
b[38222] == 38222 && 
b[38223] == 38223 && 
b[38224] == 38224 && 
b[38225] == 38225 && 
b[38226] == 38226 && 
b[38227] == 38227 && 
b[38228] == 38228 && 
b[38229] == 38229 && 
b[38230] == 38230 && 
b[38231] == 38231 && 
b[38232] == 38232 && 
b[38233] == 38233 && 
b[38234] == 38234 && 
b[38235] == 38235 && 
b[38236] == 38236 && 
b[38237] == 38237 && 
b[38238] == 38238 && 
b[38239] == 38239 && 
b[38240] == 38240 && 
b[38241] == 38241 && 
b[38242] == 38242 && 
b[38243] == 38243 && 
b[38244] == 38244 && 
b[38245] == 38245 && 
b[38246] == 38246 && 
b[38247] == 38247 && 
b[38248] == 38248 && 
b[38249] == 38249 && 
b[38250] == 38250 && 
b[38251] == 38251 && 
b[38252] == 38252 && 
b[38253] == 38253 && 
b[38254] == 38254 && 
b[38255] == 38255 && 
b[38256] == 38256 && 
b[38257] == 38257 && 
b[38258] == 38258 && 
b[38259] == 38259 && 
b[38260] == 38260 && 
b[38261] == 38261 && 
b[38262] == 38262 && 
b[38263] == 38263 && 
b[38264] == 38264 && 
b[38265] == 38265 && 
b[38266] == 38266 && 
b[38267] == 38267 && 
b[38268] == 38268 && 
b[38269] == 38269 && 
b[38270] == 38270 && 
b[38271] == 38271 && 
b[38272] == 38272 && 
b[38273] == 38273 && 
b[38274] == 38274 && 
b[38275] == 38275 && 
b[38276] == 38276 && 
b[38277] == 38277 && 
b[38278] == 38278 && 
b[38279] == 38279 && 
b[38280] == 38280 && 
b[38281] == 38281 && 
b[38282] == 38282 && 
b[38283] == 38283 && 
b[38284] == 38284 && 
b[38285] == 38285 && 
b[38286] == 38286 && 
b[38287] == 38287 && 
b[38288] == 38288 && 
b[38289] == 38289 && 
b[38290] == 38290 && 
b[38291] == 38291 && 
b[38292] == 38292 && 
b[38293] == 38293 && 
b[38294] == 38294 && 
b[38295] == 38295 && 
b[38296] == 38296 && 
b[38297] == 38297 && 
b[38298] == 38298 && 
b[38299] == 38299 && 
b[38300] == 38300 && 
b[38301] == 38301 && 
b[38302] == 38302 && 
b[38303] == 38303 && 
b[38304] == 38304 && 
b[38305] == 38305 && 
b[38306] == 38306 && 
b[38307] == 38307 && 
b[38308] == 38308 && 
b[38309] == 38309 && 
b[38310] == 38310 && 
b[38311] == 38311 && 
b[38312] == 38312 && 
b[38313] == 38313 && 
b[38314] == 38314 && 
b[38315] == 38315 && 
b[38316] == 38316 && 
b[38317] == 38317 && 
b[38318] == 38318 && 
b[38319] == 38319 && 
b[38320] == 38320 && 
b[38321] == 38321 && 
b[38322] == 38322 && 
b[38323] == 38323 && 
b[38324] == 38324 && 
b[38325] == 38325 && 
b[38326] == 38326 && 
b[38327] == 38327 && 
b[38328] == 38328 && 
b[38329] == 38329 && 
b[38330] == 38330 && 
b[38331] == 38331 && 
b[38332] == 38332 && 
b[38333] == 38333 && 
b[38334] == 38334 && 
b[38335] == 38335 && 
b[38336] == 38336 && 
b[38337] == 38337 && 
b[38338] == 38338 && 
b[38339] == 38339 && 
b[38340] == 38340 && 
b[38341] == 38341 && 
b[38342] == 38342 && 
b[38343] == 38343 && 
b[38344] == 38344 && 
b[38345] == 38345 && 
b[38346] == 38346 && 
b[38347] == 38347 && 
b[38348] == 38348 && 
b[38349] == 38349 && 
b[38350] == 38350 && 
b[38351] == 38351 && 
b[38352] == 38352 && 
b[38353] == 38353 && 
b[38354] == 38354 && 
b[38355] == 38355 && 
b[38356] == 38356 && 
b[38357] == 38357 && 
b[38358] == 38358 && 
b[38359] == 38359 && 
b[38360] == 38360 && 
b[38361] == 38361 && 
b[38362] == 38362 && 
b[38363] == 38363 && 
b[38364] == 38364 && 
b[38365] == 38365 && 
b[38366] == 38366 && 
b[38367] == 38367 && 
b[38368] == 38368 && 
b[38369] == 38369 && 
b[38370] == 38370 && 
b[38371] == 38371 && 
b[38372] == 38372 && 
b[38373] == 38373 && 
b[38374] == 38374 && 
b[38375] == 38375 && 
b[38376] == 38376 && 
b[38377] == 38377 && 
b[38378] == 38378 && 
b[38379] == 38379 && 
b[38380] == 38380 && 
b[38381] == 38381 && 
b[38382] == 38382 && 
b[38383] == 38383 && 
b[38384] == 38384 && 
b[38385] == 38385 && 
b[38386] == 38386 && 
b[38387] == 38387 && 
b[38388] == 38388 && 
b[38389] == 38389 && 
b[38390] == 38390 && 
b[38391] == 38391 && 
b[38392] == 38392 && 
b[38393] == 38393 && 
b[38394] == 38394 && 
b[38395] == 38395 && 
b[38396] == 38396 && 
b[38397] == 38397 && 
b[38398] == 38398 && 
b[38399] == 38399 && 
b[38400] == 38400 && 
b[38401] == 38401 && 
b[38402] == 38402 && 
b[38403] == 38403 && 
b[38404] == 38404 && 
b[38405] == 38405 && 
b[38406] == 38406 && 
b[38407] == 38407 && 
b[38408] == 38408 && 
b[38409] == 38409 && 
b[38410] == 38410 && 
b[38411] == 38411 && 
b[38412] == 38412 && 
b[38413] == 38413 && 
b[38414] == 38414 && 
b[38415] == 38415 && 
b[38416] == 38416 && 
b[38417] == 38417 && 
b[38418] == 38418 && 
b[38419] == 38419 && 
b[38420] == 38420 && 
b[38421] == 38421 && 
b[38422] == 38422 && 
b[38423] == 38423 && 
b[38424] == 38424 && 
b[38425] == 38425 && 
b[38426] == 38426 && 
b[38427] == 38427 && 
b[38428] == 38428 && 
b[38429] == 38429 && 
b[38430] == 38430 && 
b[38431] == 38431 && 
b[38432] == 38432 && 
b[38433] == 38433 && 
b[38434] == 38434 && 
b[38435] == 38435 && 
b[38436] == 38436 && 
b[38437] == 38437 && 
b[38438] == 38438 && 
b[38439] == 38439 && 
b[38440] == 38440 && 
b[38441] == 38441 && 
b[38442] == 38442 && 
b[38443] == 38443 && 
b[38444] == 38444 && 
b[38445] == 38445 && 
b[38446] == 38446 && 
b[38447] == 38447 && 
b[38448] == 38448 && 
b[38449] == 38449 && 
b[38450] == 38450 && 
b[38451] == 38451 && 
b[38452] == 38452 && 
b[38453] == 38453 && 
b[38454] == 38454 && 
b[38455] == 38455 && 
b[38456] == 38456 && 
b[38457] == 38457 && 
b[38458] == 38458 && 
b[38459] == 38459 && 
b[38460] == 38460 && 
b[38461] == 38461 && 
b[38462] == 38462 && 
b[38463] == 38463 && 
b[38464] == 38464 && 
b[38465] == 38465 && 
b[38466] == 38466 && 
b[38467] == 38467 && 
b[38468] == 38468 && 
b[38469] == 38469 && 
b[38470] == 38470 && 
b[38471] == 38471 && 
b[38472] == 38472 && 
b[38473] == 38473 && 
b[38474] == 38474 && 
b[38475] == 38475 && 
b[38476] == 38476 && 
b[38477] == 38477 && 
b[38478] == 38478 && 
b[38479] == 38479 && 
b[38480] == 38480 && 
b[38481] == 38481 && 
b[38482] == 38482 && 
b[38483] == 38483 && 
b[38484] == 38484 && 
b[38485] == 38485 && 
b[38486] == 38486 && 
b[38487] == 38487 && 
b[38488] == 38488 && 
b[38489] == 38489 && 
b[38490] == 38490 && 
b[38491] == 38491 && 
b[38492] == 38492 && 
b[38493] == 38493 && 
b[38494] == 38494 && 
b[38495] == 38495 && 
b[38496] == 38496 && 
b[38497] == 38497 && 
b[38498] == 38498 && 
b[38499] == 38499 && 
b[38500] == 38500 && 
b[38501] == 38501 && 
b[38502] == 38502 && 
b[38503] == 38503 && 
b[38504] == 38504 && 
b[38505] == 38505 && 
b[38506] == 38506 && 
b[38507] == 38507 && 
b[38508] == 38508 && 
b[38509] == 38509 && 
b[38510] == 38510 && 
b[38511] == 38511 && 
b[38512] == 38512 && 
b[38513] == 38513 && 
b[38514] == 38514 && 
b[38515] == 38515 && 
b[38516] == 38516 && 
b[38517] == 38517 && 
b[38518] == 38518 && 
b[38519] == 38519 && 
b[38520] == 38520 && 
b[38521] == 38521 && 
b[38522] == 38522 && 
b[38523] == 38523 && 
b[38524] == 38524 && 
b[38525] == 38525 && 
b[38526] == 38526 && 
b[38527] == 38527 && 
b[38528] == 38528 && 
b[38529] == 38529 && 
b[38530] == 38530 && 
b[38531] == 38531 && 
b[38532] == 38532 && 
b[38533] == 38533 && 
b[38534] == 38534 && 
b[38535] == 38535 && 
b[38536] == 38536 && 
b[38537] == 38537 && 
b[38538] == 38538 && 
b[38539] == 38539 && 
b[38540] == 38540 && 
b[38541] == 38541 && 
b[38542] == 38542 && 
b[38543] == 38543 && 
b[38544] == 38544 && 
b[38545] == 38545 && 
b[38546] == 38546 && 
b[38547] == 38547 && 
b[38548] == 38548 && 
b[38549] == 38549 && 
b[38550] == 38550 && 
b[38551] == 38551 && 
b[38552] == 38552 && 
b[38553] == 38553 && 
b[38554] == 38554 && 
b[38555] == 38555 && 
b[38556] == 38556 && 
b[38557] == 38557 && 
b[38558] == 38558 && 
b[38559] == 38559 && 
b[38560] == 38560 && 
b[38561] == 38561 && 
b[38562] == 38562 && 
b[38563] == 38563 && 
b[38564] == 38564 && 
b[38565] == 38565 && 
b[38566] == 38566 && 
b[38567] == 38567 && 
b[38568] == 38568 && 
b[38569] == 38569 && 
b[38570] == 38570 && 
b[38571] == 38571 && 
b[38572] == 38572 && 
b[38573] == 38573 && 
b[38574] == 38574 && 
b[38575] == 38575 && 
b[38576] == 38576 && 
b[38577] == 38577 && 
b[38578] == 38578 && 
b[38579] == 38579 && 
b[38580] == 38580 && 
b[38581] == 38581 && 
b[38582] == 38582 && 
b[38583] == 38583 && 
b[38584] == 38584 && 
b[38585] == 38585 && 
b[38586] == 38586 && 
b[38587] == 38587 && 
b[38588] == 38588 && 
b[38589] == 38589 && 
b[38590] == 38590 && 
b[38591] == 38591 && 
b[38592] == 38592 && 
b[38593] == 38593 && 
b[38594] == 38594 && 
b[38595] == 38595 && 
b[38596] == 38596 && 
b[38597] == 38597 && 
b[38598] == 38598 && 
b[38599] == 38599 && 
b[38600] == 38600 && 
b[38601] == 38601 && 
b[38602] == 38602 && 
b[38603] == 38603 && 
b[38604] == 38604 && 
b[38605] == 38605 && 
b[38606] == 38606 && 
b[38607] == 38607 && 
b[38608] == 38608 && 
b[38609] == 38609 && 
b[38610] == 38610 && 
b[38611] == 38611 && 
b[38612] == 38612 && 
b[38613] == 38613 && 
b[38614] == 38614 && 
b[38615] == 38615 && 
b[38616] == 38616 && 
b[38617] == 38617 && 
b[38618] == 38618 && 
b[38619] == 38619 && 
b[38620] == 38620 && 
b[38621] == 38621 && 
b[38622] == 38622 && 
b[38623] == 38623 && 
b[38624] == 38624 && 
b[38625] == 38625 && 
b[38626] == 38626 && 
b[38627] == 38627 && 
b[38628] == 38628 && 
b[38629] == 38629 && 
b[38630] == 38630 && 
b[38631] == 38631 && 
b[38632] == 38632 && 
b[38633] == 38633 && 
b[38634] == 38634 && 
b[38635] == 38635 && 
b[38636] == 38636 && 
b[38637] == 38637 && 
b[38638] == 38638 && 
b[38639] == 38639 && 
b[38640] == 38640 && 
b[38641] == 38641 && 
b[38642] == 38642 && 
b[38643] == 38643 && 
b[38644] == 38644 && 
b[38645] == 38645 && 
b[38646] == 38646 && 
b[38647] == 38647 && 
b[38648] == 38648 && 
b[38649] == 38649 && 
b[38650] == 38650 && 
b[38651] == 38651 && 
b[38652] == 38652 && 
b[38653] == 38653 && 
b[38654] == 38654 && 
b[38655] == 38655 && 
b[38656] == 38656 && 
b[38657] == 38657 && 
b[38658] == 38658 && 
b[38659] == 38659 && 
b[38660] == 38660 && 
b[38661] == 38661 && 
b[38662] == 38662 && 
b[38663] == 38663 && 
b[38664] == 38664 && 
b[38665] == 38665 && 
b[38666] == 38666 && 
b[38667] == 38667 && 
b[38668] == 38668 && 
b[38669] == 38669 && 
b[38670] == 38670 && 
b[38671] == 38671 && 
b[38672] == 38672 && 
b[38673] == 38673 && 
b[38674] == 38674 && 
b[38675] == 38675 && 
b[38676] == 38676 && 
b[38677] == 38677 && 
b[38678] == 38678 && 
b[38679] == 38679 && 
b[38680] == 38680 && 
b[38681] == 38681 && 
b[38682] == 38682 && 
b[38683] == 38683 && 
b[38684] == 38684 && 
b[38685] == 38685 && 
b[38686] == 38686 && 
b[38687] == 38687 && 
b[38688] == 38688 && 
b[38689] == 38689 && 
b[38690] == 38690 && 
b[38691] == 38691 && 
b[38692] == 38692 && 
b[38693] == 38693 && 
b[38694] == 38694 && 
b[38695] == 38695 && 
b[38696] == 38696 && 
b[38697] == 38697 && 
b[38698] == 38698 && 
b[38699] == 38699 && 
b[38700] == 38700 && 
b[38701] == 38701 && 
b[38702] == 38702 && 
b[38703] == 38703 && 
b[38704] == 38704 && 
b[38705] == 38705 && 
b[38706] == 38706 && 
b[38707] == 38707 && 
b[38708] == 38708 && 
b[38709] == 38709 && 
b[38710] == 38710 && 
b[38711] == 38711 && 
b[38712] == 38712 && 
b[38713] == 38713 && 
b[38714] == 38714 && 
b[38715] == 38715 && 
b[38716] == 38716 && 
b[38717] == 38717 && 
b[38718] == 38718 && 
b[38719] == 38719 && 
b[38720] == 38720 && 
b[38721] == 38721 && 
b[38722] == 38722 && 
b[38723] == 38723 && 
b[38724] == 38724 && 
b[38725] == 38725 && 
b[38726] == 38726 && 
b[38727] == 38727 && 
b[38728] == 38728 && 
b[38729] == 38729 && 
b[38730] == 38730 && 
b[38731] == 38731 && 
b[38732] == 38732 && 
b[38733] == 38733 && 
b[38734] == 38734 && 
b[38735] == 38735 && 
b[38736] == 38736 && 
b[38737] == 38737 && 
b[38738] == 38738 && 
b[38739] == 38739 && 
b[38740] == 38740 && 
b[38741] == 38741 && 
b[38742] == 38742 && 
b[38743] == 38743 && 
b[38744] == 38744 && 
b[38745] == 38745 && 
b[38746] == 38746 && 
b[38747] == 38747 && 
b[38748] == 38748 && 
b[38749] == 38749 && 
b[38750] == 38750 && 
b[38751] == 38751 && 
b[38752] == 38752 && 
b[38753] == 38753 && 
b[38754] == 38754 && 
b[38755] == 38755 && 
b[38756] == 38756 && 
b[38757] == 38757 && 
b[38758] == 38758 && 
b[38759] == 38759 && 
b[38760] == 38760 && 
b[38761] == 38761 && 
b[38762] == 38762 && 
b[38763] == 38763 && 
b[38764] == 38764 && 
b[38765] == 38765 && 
b[38766] == 38766 && 
b[38767] == 38767 && 
b[38768] == 38768 && 
b[38769] == 38769 && 
b[38770] == 38770 && 
b[38771] == 38771 && 
b[38772] == 38772 && 
b[38773] == 38773 && 
b[38774] == 38774 && 
b[38775] == 38775 && 
b[38776] == 38776 && 
b[38777] == 38777 && 
b[38778] == 38778 && 
b[38779] == 38779 && 
b[38780] == 38780 && 
b[38781] == 38781 && 
b[38782] == 38782 && 
b[38783] == 38783 && 
b[38784] == 38784 && 
b[38785] == 38785 && 
b[38786] == 38786 && 
b[38787] == 38787 && 
b[38788] == 38788 && 
b[38789] == 38789 && 
b[38790] == 38790 && 
b[38791] == 38791 && 
b[38792] == 38792 && 
b[38793] == 38793 && 
b[38794] == 38794 && 
b[38795] == 38795 && 
b[38796] == 38796 && 
b[38797] == 38797 && 
b[38798] == 38798 && 
b[38799] == 38799 && 
b[38800] == 38800 && 
b[38801] == 38801 && 
b[38802] == 38802 && 
b[38803] == 38803 && 
b[38804] == 38804 && 
b[38805] == 38805 && 
b[38806] == 38806 && 
b[38807] == 38807 && 
b[38808] == 38808 && 
b[38809] == 38809 && 
b[38810] == 38810 && 
b[38811] == 38811 && 
b[38812] == 38812 && 
b[38813] == 38813 && 
b[38814] == 38814 && 
b[38815] == 38815 && 
b[38816] == 38816 && 
b[38817] == 38817 && 
b[38818] == 38818 && 
b[38819] == 38819 && 
b[38820] == 38820 && 
b[38821] == 38821 && 
b[38822] == 38822 && 
b[38823] == 38823 && 
b[38824] == 38824 && 
b[38825] == 38825 && 
b[38826] == 38826 && 
b[38827] == 38827 && 
b[38828] == 38828 && 
b[38829] == 38829 && 
b[38830] == 38830 && 
b[38831] == 38831 && 
b[38832] == 38832 && 
b[38833] == 38833 && 
b[38834] == 38834 && 
b[38835] == 38835 && 
b[38836] == 38836 && 
b[38837] == 38837 && 
b[38838] == 38838 && 
b[38839] == 38839 && 
b[38840] == 38840 && 
b[38841] == 38841 && 
b[38842] == 38842 && 
b[38843] == 38843 && 
b[38844] == 38844 && 
b[38845] == 38845 && 
b[38846] == 38846 && 
b[38847] == 38847 && 
b[38848] == 38848 && 
b[38849] == 38849 && 
b[38850] == 38850 && 
b[38851] == 38851 && 
b[38852] == 38852 && 
b[38853] == 38853 && 
b[38854] == 38854 && 
b[38855] == 38855 && 
b[38856] == 38856 && 
b[38857] == 38857 && 
b[38858] == 38858 && 
b[38859] == 38859 && 
b[38860] == 38860 && 
b[38861] == 38861 && 
b[38862] == 38862 && 
b[38863] == 38863 && 
b[38864] == 38864 && 
b[38865] == 38865 && 
b[38866] == 38866 && 
b[38867] == 38867 && 
b[38868] == 38868 && 
b[38869] == 38869 && 
b[38870] == 38870 && 
b[38871] == 38871 && 
b[38872] == 38872 && 
b[38873] == 38873 && 
b[38874] == 38874 && 
b[38875] == 38875 && 
b[38876] == 38876 && 
b[38877] == 38877 && 
b[38878] == 38878 && 
b[38879] == 38879 && 
b[38880] == 38880 && 
b[38881] == 38881 && 
b[38882] == 38882 && 
b[38883] == 38883 && 
b[38884] == 38884 && 
b[38885] == 38885 && 
b[38886] == 38886 && 
b[38887] == 38887 && 
b[38888] == 38888 && 
b[38889] == 38889 && 
b[38890] == 38890 && 
b[38891] == 38891 && 
b[38892] == 38892 && 
b[38893] == 38893 && 
b[38894] == 38894 && 
b[38895] == 38895 && 
b[38896] == 38896 && 
b[38897] == 38897 && 
b[38898] == 38898 && 
b[38899] == 38899 && 
b[38900] == 38900 && 
b[38901] == 38901 && 
b[38902] == 38902 && 
b[38903] == 38903 && 
b[38904] == 38904 && 
b[38905] == 38905 && 
b[38906] == 38906 && 
b[38907] == 38907 && 
b[38908] == 38908 && 
b[38909] == 38909 && 
b[38910] == 38910 && 
b[38911] == 38911 && 
b[38912] == 38912 && 
b[38913] == 38913 && 
b[38914] == 38914 && 
b[38915] == 38915 && 
b[38916] == 38916 && 
b[38917] == 38917 && 
b[38918] == 38918 && 
b[38919] == 38919 && 
b[38920] == 38920 && 
b[38921] == 38921 && 
b[38922] == 38922 && 
b[38923] == 38923 && 
b[38924] == 38924 && 
b[38925] == 38925 && 
b[38926] == 38926 && 
b[38927] == 38927 && 
b[38928] == 38928 && 
b[38929] == 38929 && 
b[38930] == 38930 && 
b[38931] == 38931 && 
b[38932] == 38932 && 
b[38933] == 38933 && 
b[38934] == 38934 && 
b[38935] == 38935 && 
b[38936] == 38936 && 
b[38937] == 38937 && 
b[38938] == 38938 && 
b[38939] == 38939 && 
b[38940] == 38940 && 
b[38941] == 38941 && 
b[38942] == 38942 && 
b[38943] == 38943 && 
b[38944] == 38944 && 
b[38945] == 38945 && 
b[38946] == 38946 && 
b[38947] == 38947 && 
b[38948] == 38948 && 
b[38949] == 38949 && 
b[38950] == 38950 && 
b[38951] == 38951 && 
b[38952] == 38952 && 
b[38953] == 38953 && 
b[38954] == 38954 && 
b[38955] == 38955 && 
b[38956] == 38956 && 
b[38957] == 38957 && 
b[38958] == 38958 && 
b[38959] == 38959 && 
b[38960] == 38960 && 
b[38961] == 38961 && 
b[38962] == 38962 && 
b[38963] == 38963 && 
b[38964] == 38964 && 
b[38965] == 38965 && 
b[38966] == 38966 && 
b[38967] == 38967 && 
b[38968] == 38968 && 
b[38969] == 38969 && 
b[38970] == 38970 && 
b[38971] == 38971 && 
b[38972] == 38972 && 
b[38973] == 38973 && 
b[38974] == 38974 && 
b[38975] == 38975 && 
b[38976] == 38976 && 
b[38977] == 38977 && 
b[38978] == 38978 && 
b[38979] == 38979 && 
b[38980] == 38980 && 
b[38981] == 38981 && 
b[38982] == 38982 && 
b[38983] == 38983 && 
b[38984] == 38984 && 
b[38985] == 38985 && 
b[38986] == 38986 && 
b[38987] == 38987 && 
b[38988] == 38988 && 
b[38989] == 38989 && 
b[38990] == 38990 && 
b[38991] == 38991 && 
b[38992] == 38992 && 
b[38993] == 38993 && 
b[38994] == 38994 && 
b[38995] == 38995 && 
b[38996] == 38996 && 
b[38997] == 38997 && 
b[38998] == 38998 && 
b[38999] == 38999 && 
b[39000] == 39000 && 
b[39001] == 39001 && 
b[39002] == 39002 && 
b[39003] == 39003 && 
b[39004] == 39004 && 
b[39005] == 39005 && 
b[39006] == 39006 && 
b[39007] == 39007 && 
b[39008] == 39008 && 
b[39009] == 39009 && 
b[39010] == 39010 && 
b[39011] == 39011 && 
b[39012] == 39012 && 
b[39013] == 39013 && 
b[39014] == 39014 && 
b[39015] == 39015 && 
b[39016] == 39016 && 
b[39017] == 39017 && 
b[39018] == 39018 && 
b[39019] == 39019 && 
b[39020] == 39020 && 
b[39021] == 39021 && 
b[39022] == 39022 && 
b[39023] == 39023 && 
b[39024] == 39024 && 
b[39025] == 39025 && 
b[39026] == 39026 && 
b[39027] == 39027 && 
b[39028] == 39028 && 
b[39029] == 39029 && 
b[39030] == 39030 && 
b[39031] == 39031 && 
b[39032] == 39032 && 
b[39033] == 39033 && 
b[39034] == 39034 && 
b[39035] == 39035 && 
b[39036] == 39036 && 
b[39037] == 39037 && 
b[39038] == 39038 && 
b[39039] == 39039 && 
b[39040] == 39040 && 
b[39041] == 39041 && 
b[39042] == 39042 && 
b[39043] == 39043 && 
b[39044] == 39044 && 
b[39045] == 39045 && 
b[39046] == 39046 && 
b[39047] == 39047 && 
b[39048] == 39048 && 
b[39049] == 39049 && 
b[39050] == 39050 && 
b[39051] == 39051 && 
b[39052] == 39052 && 
b[39053] == 39053 && 
b[39054] == 39054 && 
b[39055] == 39055 && 
b[39056] == 39056 && 
b[39057] == 39057 && 
b[39058] == 39058 && 
b[39059] == 39059 && 
b[39060] == 39060 && 
b[39061] == 39061 && 
b[39062] == 39062 && 
b[39063] == 39063 && 
b[39064] == 39064 && 
b[39065] == 39065 && 
b[39066] == 39066 && 
b[39067] == 39067 && 
b[39068] == 39068 && 
b[39069] == 39069 && 
b[39070] == 39070 && 
b[39071] == 39071 && 
b[39072] == 39072 && 
b[39073] == 39073 && 
b[39074] == 39074 && 
b[39075] == 39075 && 
b[39076] == 39076 && 
b[39077] == 39077 && 
b[39078] == 39078 && 
b[39079] == 39079 && 
b[39080] == 39080 && 
b[39081] == 39081 && 
b[39082] == 39082 && 
b[39083] == 39083 && 
b[39084] == 39084 && 
b[39085] == 39085 && 
b[39086] == 39086 && 
b[39087] == 39087 && 
b[39088] == 39088 && 
b[39089] == 39089 && 
b[39090] == 39090 && 
b[39091] == 39091 && 
b[39092] == 39092 && 
b[39093] == 39093 && 
b[39094] == 39094 && 
b[39095] == 39095 && 
b[39096] == 39096 && 
b[39097] == 39097 && 
b[39098] == 39098 && 
b[39099] == 39099 && 
b[39100] == 39100 && 
b[39101] == 39101 && 
b[39102] == 39102 && 
b[39103] == 39103 && 
b[39104] == 39104 && 
b[39105] == 39105 && 
b[39106] == 39106 && 
b[39107] == 39107 && 
b[39108] == 39108 && 
b[39109] == 39109 && 
b[39110] == 39110 && 
b[39111] == 39111 && 
b[39112] == 39112 && 
b[39113] == 39113 && 
b[39114] == 39114 && 
b[39115] == 39115 && 
b[39116] == 39116 && 
b[39117] == 39117 && 
b[39118] == 39118 && 
b[39119] == 39119 && 
b[39120] == 39120 && 
b[39121] == 39121 && 
b[39122] == 39122 && 
b[39123] == 39123 && 
b[39124] == 39124 && 
b[39125] == 39125 && 
b[39126] == 39126 && 
b[39127] == 39127 && 
b[39128] == 39128 && 
b[39129] == 39129 && 
b[39130] == 39130 && 
b[39131] == 39131 && 
b[39132] == 39132 && 
b[39133] == 39133 && 
b[39134] == 39134 && 
b[39135] == 39135 && 
b[39136] == 39136 && 
b[39137] == 39137 && 
b[39138] == 39138 && 
b[39139] == 39139 && 
b[39140] == 39140 && 
b[39141] == 39141 && 
b[39142] == 39142 && 
b[39143] == 39143 && 
b[39144] == 39144 && 
b[39145] == 39145 && 
b[39146] == 39146 && 
b[39147] == 39147 && 
b[39148] == 39148 && 
b[39149] == 39149 && 
b[39150] == 39150 && 
b[39151] == 39151 && 
b[39152] == 39152 && 
b[39153] == 39153 && 
b[39154] == 39154 && 
b[39155] == 39155 && 
b[39156] == 39156 && 
b[39157] == 39157 && 
b[39158] == 39158 && 
b[39159] == 39159 && 
b[39160] == 39160 && 
b[39161] == 39161 && 
b[39162] == 39162 && 
b[39163] == 39163 && 
b[39164] == 39164 && 
b[39165] == 39165 && 
b[39166] == 39166 && 
b[39167] == 39167 && 
b[39168] == 39168 && 
b[39169] == 39169 && 
b[39170] == 39170 && 
b[39171] == 39171 && 
b[39172] == 39172 && 
b[39173] == 39173 && 
b[39174] == 39174 && 
b[39175] == 39175 && 
b[39176] == 39176 && 
b[39177] == 39177 && 
b[39178] == 39178 && 
b[39179] == 39179 && 
b[39180] == 39180 && 
b[39181] == 39181 && 
b[39182] == 39182 && 
b[39183] == 39183 && 
b[39184] == 39184 && 
b[39185] == 39185 && 
b[39186] == 39186 && 
b[39187] == 39187 && 
b[39188] == 39188 && 
b[39189] == 39189 && 
b[39190] == 39190 && 
b[39191] == 39191 && 
b[39192] == 39192 && 
b[39193] == 39193 && 
b[39194] == 39194 && 
b[39195] == 39195 && 
b[39196] == 39196 && 
b[39197] == 39197 && 
b[39198] == 39198 && 
b[39199] == 39199 && 
b[39200] == 39200 && 
b[39201] == 39201 && 
b[39202] == 39202 && 
b[39203] == 39203 && 
b[39204] == 39204 && 
b[39205] == 39205 && 
b[39206] == 39206 && 
b[39207] == 39207 && 
b[39208] == 39208 && 
b[39209] == 39209 && 
b[39210] == 39210 && 
b[39211] == 39211 && 
b[39212] == 39212 && 
b[39213] == 39213 && 
b[39214] == 39214 && 
b[39215] == 39215 && 
b[39216] == 39216 && 
b[39217] == 39217 && 
b[39218] == 39218 && 
b[39219] == 39219 && 
b[39220] == 39220 && 
b[39221] == 39221 && 
b[39222] == 39222 && 
b[39223] == 39223 && 
b[39224] == 39224 && 
b[39225] == 39225 && 
b[39226] == 39226 && 
b[39227] == 39227 && 
b[39228] == 39228 && 
b[39229] == 39229 && 
b[39230] == 39230 && 
b[39231] == 39231 && 
b[39232] == 39232 && 
b[39233] == 39233 && 
b[39234] == 39234 && 
b[39235] == 39235 && 
b[39236] == 39236 && 
b[39237] == 39237 && 
b[39238] == 39238 && 
b[39239] == 39239 && 
b[39240] == 39240 && 
b[39241] == 39241 && 
b[39242] == 39242 && 
b[39243] == 39243 && 
b[39244] == 39244 && 
b[39245] == 39245 && 
b[39246] == 39246 && 
b[39247] == 39247 && 
b[39248] == 39248 && 
b[39249] == 39249 && 
b[39250] == 39250 && 
b[39251] == 39251 && 
b[39252] == 39252 && 
b[39253] == 39253 && 
b[39254] == 39254 && 
b[39255] == 39255 && 
b[39256] == 39256 && 
b[39257] == 39257 && 
b[39258] == 39258 && 
b[39259] == 39259 && 
b[39260] == 39260 && 
b[39261] == 39261 && 
b[39262] == 39262 && 
b[39263] == 39263 && 
b[39264] == 39264 && 
b[39265] == 39265 && 
b[39266] == 39266 && 
b[39267] == 39267 && 
b[39268] == 39268 && 
b[39269] == 39269 && 
b[39270] == 39270 && 
b[39271] == 39271 && 
b[39272] == 39272 && 
b[39273] == 39273 && 
b[39274] == 39274 && 
b[39275] == 39275 && 
b[39276] == 39276 && 
b[39277] == 39277 && 
b[39278] == 39278 && 
b[39279] == 39279 && 
b[39280] == 39280 && 
b[39281] == 39281 && 
b[39282] == 39282 && 
b[39283] == 39283 && 
b[39284] == 39284 && 
b[39285] == 39285 && 
b[39286] == 39286 && 
b[39287] == 39287 && 
b[39288] == 39288 && 
b[39289] == 39289 && 
b[39290] == 39290 && 
b[39291] == 39291 && 
b[39292] == 39292 && 
b[39293] == 39293 && 
b[39294] == 39294 && 
b[39295] == 39295 && 
b[39296] == 39296 && 
b[39297] == 39297 && 
b[39298] == 39298 && 
b[39299] == 39299 && 
b[39300] == 39300 && 
b[39301] == 39301 && 
b[39302] == 39302 && 
b[39303] == 39303 && 
b[39304] == 39304 && 
b[39305] == 39305 && 
b[39306] == 39306 && 
b[39307] == 39307 && 
b[39308] == 39308 && 
b[39309] == 39309 && 
b[39310] == 39310 && 
b[39311] == 39311 && 
b[39312] == 39312 && 
b[39313] == 39313 && 
b[39314] == 39314 && 
b[39315] == 39315 && 
b[39316] == 39316 && 
b[39317] == 39317 && 
b[39318] == 39318 && 
b[39319] == 39319 && 
b[39320] == 39320 && 
b[39321] == 39321 && 
b[39322] == 39322 && 
b[39323] == 39323 && 
b[39324] == 39324 && 
b[39325] == 39325 && 
b[39326] == 39326 && 
b[39327] == 39327 && 
b[39328] == 39328 && 
b[39329] == 39329 && 
b[39330] == 39330 && 
b[39331] == 39331 && 
b[39332] == 39332 && 
b[39333] == 39333 && 
b[39334] == 39334 && 
b[39335] == 39335 && 
b[39336] == 39336 && 
b[39337] == 39337 && 
b[39338] == 39338 && 
b[39339] == 39339 && 
b[39340] == 39340 && 
b[39341] == 39341 && 
b[39342] == 39342 && 
b[39343] == 39343 && 
b[39344] == 39344 && 
b[39345] == 39345 && 
b[39346] == 39346 && 
b[39347] == 39347 && 
b[39348] == 39348 && 
b[39349] == 39349 && 
b[39350] == 39350 && 
b[39351] == 39351 && 
b[39352] == 39352 && 
b[39353] == 39353 && 
b[39354] == 39354 && 
b[39355] == 39355 && 
b[39356] == 39356 && 
b[39357] == 39357 && 
b[39358] == 39358 && 
b[39359] == 39359 && 
b[39360] == 39360 && 
b[39361] == 39361 && 
b[39362] == 39362 && 
b[39363] == 39363 && 
b[39364] == 39364 && 
b[39365] == 39365 && 
b[39366] == 39366 && 
b[39367] == 39367 && 
b[39368] == 39368 && 
b[39369] == 39369 && 
b[39370] == 39370 && 
b[39371] == 39371 && 
b[39372] == 39372 && 
b[39373] == 39373 && 
b[39374] == 39374 && 
b[39375] == 39375 && 
b[39376] == 39376 && 
b[39377] == 39377 && 
b[39378] == 39378 && 
b[39379] == 39379 && 
b[39380] == 39380 && 
b[39381] == 39381 && 
b[39382] == 39382 && 
b[39383] == 39383 && 
b[39384] == 39384 && 
b[39385] == 39385 && 
b[39386] == 39386 && 
b[39387] == 39387 && 
b[39388] == 39388 && 
b[39389] == 39389 && 
b[39390] == 39390 && 
b[39391] == 39391 && 
b[39392] == 39392 && 
b[39393] == 39393 && 
b[39394] == 39394 && 
b[39395] == 39395 && 
b[39396] == 39396 && 
b[39397] == 39397 && 
b[39398] == 39398 && 
b[39399] == 39399 && 
b[39400] == 39400 && 
b[39401] == 39401 && 
b[39402] == 39402 && 
b[39403] == 39403 && 
b[39404] == 39404 && 
b[39405] == 39405 && 
b[39406] == 39406 && 
b[39407] == 39407 && 
b[39408] == 39408 && 
b[39409] == 39409 && 
b[39410] == 39410 && 
b[39411] == 39411 && 
b[39412] == 39412 && 
b[39413] == 39413 && 
b[39414] == 39414 && 
b[39415] == 39415 && 
b[39416] == 39416 && 
b[39417] == 39417 && 
b[39418] == 39418 && 
b[39419] == 39419 && 
b[39420] == 39420 && 
b[39421] == 39421 && 
b[39422] == 39422 && 
b[39423] == 39423 && 
b[39424] == 39424 && 
b[39425] == 39425 && 
b[39426] == 39426 && 
b[39427] == 39427 && 
b[39428] == 39428 && 
b[39429] == 39429 && 
b[39430] == 39430 && 
b[39431] == 39431 && 
b[39432] == 39432 && 
b[39433] == 39433 && 
b[39434] == 39434 && 
b[39435] == 39435 && 
b[39436] == 39436 && 
b[39437] == 39437 && 
b[39438] == 39438 && 
b[39439] == 39439 && 
b[39440] == 39440 && 
b[39441] == 39441 && 
b[39442] == 39442 && 
b[39443] == 39443 && 
b[39444] == 39444 && 
b[39445] == 39445 && 
b[39446] == 39446 && 
b[39447] == 39447 && 
b[39448] == 39448 && 
b[39449] == 39449 && 
b[39450] == 39450 && 
b[39451] == 39451 && 
b[39452] == 39452 && 
b[39453] == 39453 && 
b[39454] == 39454 && 
b[39455] == 39455 && 
b[39456] == 39456 && 
b[39457] == 39457 && 
b[39458] == 39458 && 
b[39459] == 39459 && 
b[39460] == 39460 && 
b[39461] == 39461 && 
b[39462] == 39462 && 
b[39463] == 39463 && 
b[39464] == 39464 && 
b[39465] == 39465 && 
b[39466] == 39466 && 
b[39467] == 39467 && 
b[39468] == 39468 && 
b[39469] == 39469 && 
b[39470] == 39470 && 
b[39471] == 39471 && 
b[39472] == 39472 && 
b[39473] == 39473 && 
b[39474] == 39474 && 
b[39475] == 39475 && 
b[39476] == 39476 && 
b[39477] == 39477 && 
b[39478] == 39478 && 
b[39479] == 39479 && 
b[39480] == 39480 && 
b[39481] == 39481 && 
b[39482] == 39482 && 
b[39483] == 39483 && 
b[39484] == 39484 && 
b[39485] == 39485 && 
b[39486] == 39486 && 
b[39487] == 39487 && 
b[39488] == 39488 && 
b[39489] == 39489 && 
b[39490] == 39490 && 
b[39491] == 39491 && 
b[39492] == 39492 && 
b[39493] == 39493 && 
b[39494] == 39494 && 
b[39495] == 39495 && 
b[39496] == 39496 && 
b[39497] == 39497 && 
b[39498] == 39498 && 
b[39499] == 39499 && 
b[39500] == 39500 && 
b[39501] == 39501 && 
b[39502] == 39502 && 
b[39503] == 39503 && 
b[39504] == 39504 && 
b[39505] == 39505 && 
b[39506] == 39506 && 
b[39507] == 39507 && 
b[39508] == 39508 && 
b[39509] == 39509 && 
b[39510] == 39510 && 
b[39511] == 39511 && 
b[39512] == 39512 && 
b[39513] == 39513 && 
b[39514] == 39514 && 
b[39515] == 39515 && 
b[39516] == 39516 && 
b[39517] == 39517 && 
b[39518] == 39518 && 
b[39519] == 39519 && 
b[39520] == 39520 && 
b[39521] == 39521 && 
b[39522] == 39522 && 
b[39523] == 39523 && 
b[39524] == 39524 && 
b[39525] == 39525 && 
b[39526] == 39526 && 
b[39527] == 39527 && 
b[39528] == 39528 && 
b[39529] == 39529 && 
b[39530] == 39530 && 
b[39531] == 39531 && 
b[39532] == 39532 && 
b[39533] == 39533 && 
b[39534] == 39534 && 
b[39535] == 39535 && 
b[39536] == 39536 && 
b[39537] == 39537 && 
b[39538] == 39538 && 
b[39539] == 39539 && 
b[39540] == 39540 && 
b[39541] == 39541 && 
b[39542] == 39542 && 
b[39543] == 39543 && 
b[39544] == 39544 && 
b[39545] == 39545 && 
b[39546] == 39546 && 
b[39547] == 39547 && 
b[39548] == 39548 && 
b[39549] == 39549 && 
b[39550] == 39550 && 
b[39551] == 39551 && 
b[39552] == 39552 && 
b[39553] == 39553 && 
b[39554] == 39554 && 
b[39555] == 39555 && 
b[39556] == 39556 && 
b[39557] == 39557 && 
b[39558] == 39558 && 
b[39559] == 39559 && 
b[39560] == 39560 && 
b[39561] == 39561 && 
b[39562] == 39562 && 
b[39563] == 39563 && 
b[39564] == 39564 && 
b[39565] == 39565 && 
b[39566] == 39566 && 
b[39567] == 39567 && 
b[39568] == 39568 && 
b[39569] == 39569 && 
b[39570] == 39570 && 
b[39571] == 39571 && 
b[39572] == 39572 && 
b[39573] == 39573 && 
b[39574] == 39574 && 
b[39575] == 39575 && 
b[39576] == 39576 && 
b[39577] == 39577 && 
b[39578] == 39578 && 
b[39579] == 39579 && 
b[39580] == 39580 && 
b[39581] == 39581 && 
b[39582] == 39582 && 
b[39583] == 39583 && 
b[39584] == 39584 && 
b[39585] == 39585 && 
b[39586] == 39586 && 
b[39587] == 39587 && 
b[39588] == 39588 && 
b[39589] == 39589 && 
b[39590] == 39590 && 
b[39591] == 39591 && 
b[39592] == 39592 && 
b[39593] == 39593 && 
b[39594] == 39594 && 
b[39595] == 39595 && 
b[39596] == 39596 && 
b[39597] == 39597 && 
b[39598] == 39598 && 
b[39599] == 39599 && 
b[39600] == 39600 && 
b[39601] == 39601 && 
b[39602] == 39602 && 
b[39603] == 39603 && 
b[39604] == 39604 && 
b[39605] == 39605 && 
b[39606] == 39606 && 
b[39607] == 39607 && 
b[39608] == 39608 && 
b[39609] == 39609 && 
b[39610] == 39610 && 
b[39611] == 39611 && 
b[39612] == 39612 && 
b[39613] == 39613 && 
b[39614] == 39614 && 
b[39615] == 39615 && 
b[39616] == 39616 && 
b[39617] == 39617 && 
b[39618] == 39618 && 
b[39619] == 39619 && 
b[39620] == 39620 && 
b[39621] == 39621 && 
b[39622] == 39622 && 
b[39623] == 39623 && 
b[39624] == 39624 && 
b[39625] == 39625 && 
b[39626] == 39626 && 
b[39627] == 39627 && 
b[39628] == 39628 && 
b[39629] == 39629 && 
b[39630] == 39630 && 
b[39631] == 39631 && 
b[39632] == 39632 && 
b[39633] == 39633 && 
b[39634] == 39634 && 
b[39635] == 39635 && 
b[39636] == 39636 && 
b[39637] == 39637 && 
b[39638] == 39638 && 
b[39639] == 39639 && 
b[39640] == 39640 && 
b[39641] == 39641 && 
b[39642] == 39642 && 
b[39643] == 39643 && 
b[39644] == 39644 && 
b[39645] == 39645 && 
b[39646] == 39646 && 
b[39647] == 39647 && 
b[39648] == 39648 && 
b[39649] == 39649 && 
b[39650] == 39650 && 
b[39651] == 39651 && 
b[39652] == 39652 && 
b[39653] == 39653 && 
b[39654] == 39654 && 
b[39655] == 39655 && 
b[39656] == 39656 && 
b[39657] == 39657 && 
b[39658] == 39658 && 
b[39659] == 39659 && 
b[39660] == 39660 && 
b[39661] == 39661 && 
b[39662] == 39662 && 
b[39663] == 39663 && 
b[39664] == 39664 && 
b[39665] == 39665 && 
b[39666] == 39666 && 
b[39667] == 39667 && 
b[39668] == 39668 && 
b[39669] == 39669 && 
b[39670] == 39670 && 
b[39671] == 39671 && 
b[39672] == 39672 && 
b[39673] == 39673 && 
b[39674] == 39674 && 
b[39675] == 39675 && 
b[39676] == 39676 && 
b[39677] == 39677 && 
b[39678] == 39678 && 
b[39679] == 39679 && 
b[39680] == 39680 && 
b[39681] == 39681 && 
b[39682] == 39682 && 
b[39683] == 39683 && 
b[39684] == 39684 && 
b[39685] == 39685 && 
b[39686] == 39686 && 
b[39687] == 39687 && 
b[39688] == 39688 && 
b[39689] == 39689 && 
b[39690] == 39690 && 
b[39691] == 39691 && 
b[39692] == 39692 && 
b[39693] == 39693 && 
b[39694] == 39694 && 
b[39695] == 39695 && 
b[39696] == 39696 && 
b[39697] == 39697 && 
b[39698] == 39698 && 
b[39699] == 39699 && 
b[39700] == 39700 && 
b[39701] == 39701 && 
b[39702] == 39702 && 
b[39703] == 39703 && 
b[39704] == 39704 && 
b[39705] == 39705 && 
b[39706] == 39706 && 
b[39707] == 39707 && 
b[39708] == 39708 && 
b[39709] == 39709 && 
b[39710] == 39710 && 
b[39711] == 39711 && 
b[39712] == 39712 && 
b[39713] == 39713 && 
b[39714] == 39714 && 
b[39715] == 39715 && 
b[39716] == 39716 && 
b[39717] == 39717 && 
b[39718] == 39718 && 
b[39719] == 39719 && 
b[39720] == 39720 && 
b[39721] == 39721 && 
b[39722] == 39722 && 
b[39723] == 39723 && 
b[39724] == 39724 && 
b[39725] == 39725 && 
b[39726] == 39726 && 
b[39727] == 39727 && 
b[39728] == 39728 && 
b[39729] == 39729 && 
b[39730] == 39730 && 
b[39731] == 39731 && 
b[39732] == 39732 && 
b[39733] == 39733 && 
b[39734] == 39734 && 
b[39735] == 39735 && 
b[39736] == 39736 && 
b[39737] == 39737 && 
b[39738] == 39738 && 
b[39739] == 39739 && 
b[39740] == 39740 && 
b[39741] == 39741 && 
b[39742] == 39742 && 
b[39743] == 39743 && 
b[39744] == 39744 && 
b[39745] == 39745 && 
b[39746] == 39746 && 
b[39747] == 39747 && 
b[39748] == 39748 && 
b[39749] == 39749 && 
b[39750] == 39750 && 
b[39751] == 39751 && 
b[39752] == 39752 && 
b[39753] == 39753 && 
b[39754] == 39754 && 
b[39755] == 39755 && 
b[39756] == 39756 && 
b[39757] == 39757 && 
b[39758] == 39758 && 
b[39759] == 39759 && 
b[39760] == 39760 && 
b[39761] == 39761 && 
b[39762] == 39762 && 
b[39763] == 39763 && 
b[39764] == 39764 && 
b[39765] == 39765 && 
b[39766] == 39766 && 
b[39767] == 39767 && 
b[39768] == 39768 && 
b[39769] == 39769 && 
b[39770] == 39770 && 
b[39771] == 39771 && 
b[39772] == 39772 && 
b[39773] == 39773 && 
b[39774] == 39774 && 
b[39775] == 39775 && 
b[39776] == 39776 && 
b[39777] == 39777 && 
b[39778] == 39778 && 
b[39779] == 39779 && 
b[39780] == 39780 && 
b[39781] == 39781 && 
b[39782] == 39782 && 
b[39783] == 39783 && 
b[39784] == 39784 && 
b[39785] == 39785 && 
b[39786] == 39786 && 
b[39787] == 39787 && 
b[39788] == 39788 && 
b[39789] == 39789 && 
b[39790] == 39790 && 
b[39791] == 39791 && 
b[39792] == 39792 && 
b[39793] == 39793 && 
b[39794] == 39794 && 
b[39795] == 39795 && 
b[39796] == 39796 && 
b[39797] == 39797 && 
b[39798] == 39798 && 
b[39799] == 39799 && 
b[39800] == 39800 && 
b[39801] == 39801 && 
b[39802] == 39802 && 
b[39803] == 39803 && 
b[39804] == 39804 && 
b[39805] == 39805 && 
b[39806] == 39806 && 
b[39807] == 39807 && 
b[39808] == 39808 && 
b[39809] == 39809 && 
b[39810] == 39810 && 
b[39811] == 39811 && 
b[39812] == 39812 && 
b[39813] == 39813 && 
b[39814] == 39814 && 
b[39815] == 39815 && 
b[39816] == 39816 && 
b[39817] == 39817 && 
b[39818] == 39818 && 
b[39819] == 39819 && 
b[39820] == 39820 && 
b[39821] == 39821 && 
b[39822] == 39822 && 
b[39823] == 39823 && 
b[39824] == 39824 && 
b[39825] == 39825 && 
b[39826] == 39826 && 
b[39827] == 39827 && 
b[39828] == 39828 && 
b[39829] == 39829 && 
b[39830] == 39830 && 
b[39831] == 39831 && 
b[39832] == 39832 && 
b[39833] == 39833 && 
b[39834] == 39834 && 
b[39835] == 39835 && 
b[39836] == 39836 && 
b[39837] == 39837 && 
b[39838] == 39838 && 
b[39839] == 39839 && 
b[39840] == 39840 && 
b[39841] == 39841 && 
b[39842] == 39842 && 
b[39843] == 39843 && 
b[39844] == 39844 && 
b[39845] == 39845 && 
b[39846] == 39846 && 
b[39847] == 39847 && 
b[39848] == 39848 && 
b[39849] == 39849 && 
b[39850] == 39850 && 
b[39851] == 39851 && 
b[39852] == 39852 && 
b[39853] == 39853 && 
b[39854] == 39854 && 
b[39855] == 39855 && 
b[39856] == 39856 && 
b[39857] == 39857 && 
b[39858] == 39858 && 
b[39859] == 39859 && 
b[39860] == 39860 && 
b[39861] == 39861 && 
b[39862] == 39862 && 
b[39863] == 39863 && 
b[39864] == 39864 && 
b[39865] == 39865 && 
b[39866] == 39866 && 
b[39867] == 39867 && 
b[39868] == 39868 && 
b[39869] == 39869 && 
b[39870] == 39870 && 
b[39871] == 39871 && 
b[39872] == 39872 && 
b[39873] == 39873 && 
b[39874] == 39874 && 
b[39875] == 39875 && 
b[39876] == 39876 && 
b[39877] == 39877 && 
b[39878] == 39878 && 
b[39879] == 39879 && 
b[39880] == 39880 && 
b[39881] == 39881 && 
b[39882] == 39882 && 
b[39883] == 39883 && 
b[39884] == 39884 && 
b[39885] == 39885 && 
b[39886] == 39886 && 
b[39887] == 39887 && 
b[39888] == 39888 && 
b[39889] == 39889 && 
b[39890] == 39890 && 
b[39891] == 39891 && 
b[39892] == 39892 && 
b[39893] == 39893 && 
b[39894] == 39894 && 
b[39895] == 39895 && 
b[39896] == 39896 && 
b[39897] == 39897 && 
b[39898] == 39898 && 
b[39899] == 39899 && 
b[39900] == 39900 && 
b[39901] == 39901 && 
b[39902] == 39902 && 
b[39903] == 39903 && 
b[39904] == 39904 && 
b[39905] == 39905 && 
b[39906] == 39906 && 
b[39907] == 39907 && 
b[39908] == 39908 && 
b[39909] == 39909 && 
b[39910] == 39910 && 
b[39911] == 39911 && 
b[39912] == 39912 && 
b[39913] == 39913 && 
b[39914] == 39914 && 
b[39915] == 39915 && 
b[39916] == 39916 && 
b[39917] == 39917 && 
b[39918] == 39918 && 
b[39919] == 39919 && 
b[39920] == 39920 && 
b[39921] == 39921 && 
b[39922] == 39922 && 
b[39923] == 39923 && 
b[39924] == 39924 && 
b[39925] == 39925 && 
b[39926] == 39926 && 
b[39927] == 39927 && 
b[39928] == 39928 && 
b[39929] == 39929 && 
b[39930] == 39930 && 
b[39931] == 39931 && 
b[39932] == 39932 && 
b[39933] == 39933 && 
b[39934] == 39934 && 
b[39935] == 39935 && 
b[39936] == 39936 && 
b[39937] == 39937 && 
b[39938] == 39938 && 
b[39939] == 39939 && 
b[39940] == 39940 && 
b[39941] == 39941 && 
b[39942] == 39942 && 
b[39943] == 39943 && 
b[39944] == 39944 && 
b[39945] == 39945 && 
b[39946] == 39946 && 
b[39947] == 39947 && 
b[39948] == 39948 && 
b[39949] == 39949 && 
b[39950] == 39950 && 
b[39951] == 39951 && 
b[39952] == 39952 && 
b[39953] == 39953 && 
b[39954] == 39954 && 
b[39955] == 39955 && 
b[39956] == 39956 && 
b[39957] == 39957 && 
b[39958] == 39958 && 
b[39959] == 39959 && 
b[39960] == 39960 && 
b[39961] == 39961 && 
b[39962] == 39962 && 
b[39963] == 39963 && 
b[39964] == 39964 && 
b[39965] == 39965 && 
b[39966] == 39966 && 
b[39967] == 39967 && 
b[39968] == 39968 && 
b[39969] == 39969 && 
b[39970] == 39970 && 
b[39971] == 39971 && 
b[39972] == 39972 && 
b[39973] == 39973 && 
b[39974] == 39974 && 
b[39975] == 39975 && 
b[39976] == 39976 && 
b[39977] == 39977 && 
b[39978] == 39978 && 
b[39979] == 39979 && 
b[39980] == 39980 && 
b[39981] == 39981 && 
b[39982] == 39982 && 
b[39983] == 39983 && 
b[39984] == 39984 && 
b[39985] == 39985 && 
b[39986] == 39986 && 
b[39987] == 39987 && 
b[39988] == 39988 && 
b[39989] == 39989 && 
b[39990] == 39990 && 
b[39991] == 39991 && 
b[39992] == 39992 && 
b[39993] == 39993 && 
b[39994] == 39994 && 
b[39995] == 39995 && 
b[39996] == 39996 && 
b[39997] == 39997 && 
b[39998] == 39998 && 
b[39999] == 39999 && 
b[40000] == 40000 && 
b[40001] == 40001 && 
b[40002] == 40002 && 
b[40003] == 40003 && 
b[40004] == 40004 && 
b[40005] == 40005 && 
b[40006] == 40006 && 
b[40007] == 40007 && 
b[40008] == 40008 && 
b[40009] == 40009 && 
b[40010] == 40010 && 
b[40011] == 40011 && 
b[40012] == 40012 && 
b[40013] == 40013 && 
b[40014] == 40014 && 
b[40015] == 40015 && 
b[40016] == 40016 && 
b[40017] == 40017 && 
b[40018] == 40018 && 
b[40019] == 40019 && 
b[40020] == 40020 && 
b[40021] == 40021 && 
b[40022] == 40022 && 
b[40023] == 40023 && 
b[40024] == 40024 && 
b[40025] == 40025 && 
b[40026] == 40026 && 
b[40027] == 40027 && 
b[40028] == 40028 && 
b[40029] == 40029 && 
b[40030] == 40030 && 
b[40031] == 40031 && 
b[40032] == 40032 && 
b[40033] == 40033 && 
b[40034] == 40034 && 
b[40035] == 40035 && 
b[40036] == 40036 && 
b[40037] == 40037 && 
b[40038] == 40038 && 
b[40039] == 40039 && 
b[40040] == 40040 && 
b[40041] == 40041 && 
b[40042] == 40042 && 
b[40043] == 40043 && 
b[40044] == 40044 && 
b[40045] == 40045 && 
b[40046] == 40046 && 
b[40047] == 40047 && 
b[40048] == 40048 && 
b[40049] == 40049 && 
b[40050] == 40050 && 
b[40051] == 40051 && 
b[40052] == 40052 && 
b[40053] == 40053 && 
b[40054] == 40054 && 
b[40055] == 40055 && 
b[40056] == 40056 && 
b[40057] == 40057 && 
b[40058] == 40058 && 
b[40059] == 40059 && 
b[40060] == 40060 && 
b[40061] == 40061 && 
b[40062] == 40062 && 
b[40063] == 40063 && 
b[40064] == 40064 && 
b[40065] == 40065 && 
b[40066] == 40066 && 
b[40067] == 40067 && 
b[40068] == 40068 && 
b[40069] == 40069 && 
b[40070] == 40070 && 
b[40071] == 40071 && 
b[40072] == 40072 && 
b[40073] == 40073 && 
b[40074] == 40074 && 
b[40075] == 40075 && 
b[40076] == 40076 && 
b[40077] == 40077 && 
b[40078] == 40078 && 
b[40079] == 40079 && 
b[40080] == 40080 && 
b[40081] == 40081 && 
b[40082] == 40082 && 
b[40083] == 40083 && 
b[40084] == 40084 && 
b[40085] == 40085 && 
b[40086] == 40086 && 
b[40087] == 40087 && 
b[40088] == 40088 && 
b[40089] == 40089 && 
b[40090] == 40090 && 
b[40091] == 40091 && 
b[40092] == 40092 && 
b[40093] == 40093 && 
b[40094] == 40094 && 
b[40095] == 40095 && 
b[40096] == 40096 && 
b[40097] == 40097 && 
b[40098] == 40098 && 
b[40099] == 40099 && 
b[40100] == 40100 && 
b[40101] == 40101 && 
b[40102] == 40102 && 
b[40103] == 40103 && 
b[40104] == 40104 && 
b[40105] == 40105 && 
b[40106] == 40106 && 
b[40107] == 40107 && 
b[40108] == 40108 && 
b[40109] == 40109 && 
b[40110] == 40110 && 
b[40111] == 40111 && 
b[40112] == 40112 && 
b[40113] == 40113 && 
b[40114] == 40114 && 
b[40115] == 40115 && 
b[40116] == 40116 && 
b[40117] == 40117 && 
b[40118] == 40118 && 
b[40119] == 40119 && 
b[40120] == 40120 && 
b[40121] == 40121 && 
b[40122] == 40122 && 
b[40123] == 40123 && 
b[40124] == 40124 && 
b[40125] == 40125 && 
b[40126] == 40126 && 
b[40127] == 40127 && 
b[40128] == 40128 && 
b[40129] == 40129 && 
b[40130] == 40130 && 
b[40131] == 40131 && 
b[40132] == 40132 && 
b[40133] == 40133 && 
b[40134] == 40134 && 
b[40135] == 40135 && 
b[40136] == 40136 && 
b[40137] == 40137 && 
b[40138] == 40138 && 
b[40139] == 40139 && 
b[40140] == 40140 && 
b[40141] == 40141 && 
b[40142] == 40142 && 
b[40143] == 40143 && 
b[40144] == 40144 && 
b[40145] == 40145 && 
b[40146] == 40146 && 
b[40147] == 40147 && 
b[40148] == 40148 && 
b[40149] == 40149 && 
b[40150] == 40150 && 
b[40151] == 40151 && 
b[40152] == 40152 && 
b[40153] == 40153 && 
b[40154] == 40154 && 
b[40155] == 40155 && 
b[40156] == 40156 && 
b[40157] == 40157 && 
b[40158] == 40158 && 
b[40159] == 40159 && 
b[40160] == 40160 && 
b[40161] == 40161 && 
b[40162] == 40162 && 
b[40163] == 40163 && 
b[40164] == 40164 && 
b[40165] == 40165 && 
b[40166] == 40166 && 
b[40167] == 40167 && 
b[40168] == 40168 && 
b[40169] == 40169 && 
b[40170] == 40170 && 
b[40171] == 40171 && 
b[40172] == 40172 && 
b[40173] == 40173 && 
b[40174] == 40174 && 
b[40175] == 40175 && 
b[40176] == 40176 && 
b[40177] == 40177 && 
b[40178] == 40178 && 
b[40179] == 40179 && 
b[40180] == 40180 && 
b[40181] == 40181 && 
b[40182] == 40182 && 
b[40183] == 40183 && 
b[40184] == 40184 && 
b[40185] == 40185 && 
b[40186] == 40186 && 
b[40187] == 40187 && 
b[40188] == 40188 && 
b[40189] == 40189 && 
b[40190] == 40190 && 
b[40191] == 40191 && 
b[40192] == 40192 && 
b[40193] == 40193 && 
b[40194] == 40194 && 
b[40195] == 40195 && 
b[40196] == 40196 && 
b[40197] == 40197 && 
b[40198] == 40198 && 
b[40199] == 40199 && 
b[40200] == 40200 && 
b[40201] == 40201 && 
b[40202] == 40202 && 
b[40203] == 40203 && 
b[40204] == 40204 && 
b[40205] == 40205 && 
b[40206] == 40206 && 
b[40207] == 40207 && 
b[40208] == 40208 && 
b[40209] == 40209 && 
b[40210] == 40210 && 
b[40211] == 40211 && 
b[40212] == 40212 && 
b[40213] == 40213 && 
b[40214] == 40214 && 
b[40215] == 40215 && 
b[40216] == 40216 && 
b[40217] == 40217 && 
b[40218] == 40218 && 
b[40219] == 40219 && 
b[40220] == 40220 && 
b[40221] == 40221 && 
b[40222] == 40222 && 
b[40223] == 40223 && 
b[40224] == 40224 && 
b[40225] == 40225 && 
b[40226] == 40226 && 
b[40227] == 40227 && 
b[40228] == 40228 && 
b[40229] == 40229 && 
b[40230] == 40230 && 
b[40231] == 40231 && 
b[40232] == 40232 && 
b[40233] == 40233 && 
b[40234] == 40234 && 
b[40235] == 40235 && 
b[40236] == 40236 && 
b[40237] == 40237 && 
b[40238] == 40238 && 
b[40239] == 40239 && 
b[40240] == 40240 && 
b[40241] == 40241 && 
b[40242] == 40242 && 
b[40243] == 40243 && 
b[40244] == 40244 && 
b[40245] == 40245 && 
b[40246] == 40246 && 
b[40247] == 40247 && 
b[40248] == 40248 && 
b[40249] == 40249 && 
b[40250] == 40250 && 
b[40251] == 40251 && 
b[40252] == 40252 && 
b[40253] == 40253 && 
b[40254] == 40254 && 
b[40255] == 40255 && 
b[40256] == 40256 && 
b[40257] == 40257 && 
b[40258] == 40258 && 
b[40259] == 40259 && 
b[40260] == 40260 && 
b[40261] == 40261 && 
b[40262] == 40262 && 
b[40263] == 40263 && 
b[40264] == 40264 && 
b[40265] == 40265 && 
b[40266] == 40266 && 
b[40267] == 40267 && 
b[40268] == 40268 && 
b[40269] == 40269 && 
b[40270] == 40270 && 
b[40271] == 40271 && 
b[40272] == 40272 && 
b[40273] == 40273 && 
b[40274] == 40274 && 
b[40275] == 40275 && 
b[40276] == 40276 && 
b[40277] == 40277 && 
b[40278] == 40278 && 
b[40279] == 40279 && 
b[40280] == 40280 && 
b[40281] == 40281 && 
b[40282] == 40282 && 
b[40283] == 40283 && 
b[40284] == 40284 && 
b[40285] == 40285 && 
b[40286] == 40286 && 
b[40287] == 40287 && 
b[40288] == 40288 && 
b[40289] == 40289 && 
b[40290] == 40290 && 
b[40291] == 40291 && 
b[40292] == 40292 && 
b[40293] == 40293 && 
b[40294] == 40294 && 
b[40295] == 40295 && 
b[40296] == 40296 && 
b[40297] == 40297 && 
b[40298] == 40298 && 
b[40299] == 40299 && 
b[40300] == 40300 && 
b[40301] == 40301 && 
b[40302] == 40302 && 
b[40303] == 40303 && 
b[40304] == 40304 && 
b[40305] == 40305 && 
b[40306] == 40306 && 
b[40307] == 40307 && 
b[40308] == 40308 && 
b[40309] == 40309 && 
b[40310] == 40310 && 
b[40311] == 40311 && 
b[40312] == 40312 && 
b[40313] == 40313 && 
b[40314] == 40314 && 
b[40315] == 40315 && 
b[40316] == 40316 && 
b[40317] == 40317 && 
b[40318] == 40318 && 
b[40319] == 40319 && 
b[40320] == 40320 && 
b[40321] == 40321 && 
b[40322] == 40322 && 
b[40323] == 40323 && 
b[40324] == 40324 && 
b[40325] == 40325 && 
b[40326] == 40326 && 
b[40327] == 40327 && 
b[40328] == 40328 && 
b[40329] == 40329 && 
b[40330] == 40330 && 
b[40331] == 40331 && 
b[40332] == 40332 && 
b[40333] == 40333 && 
b[40334] == 40334 && 
b[40335] == 40335 && 
b[40336] == 40336 && 
b[40337] == 40337 && 
b[40338] == 40338 && 
b[40339] == 40339 && 
b[40340] == 40340 && 
b[40341] == 40341 && 
b[40342] == 40342 && 
b[40343] == 40343 && 
b[40344] == 40344 && 
b[40345] == 40345 && 
b[40346] == 40346 && 
b[40347] == 40347 && 
b[40348] == 40348 && 
b[40349] == 40349 && 
b[40350] == 40350 && 
b[40351] == 40351 && 
b[40352] == 40352 && 
b[40353] == 40353 && 
b[40354] == 40354 && 
b[40355] == 40355 && 
b[40356] == 40356 && 
b[40357] == 40357 && 
b[40358] == 40358 && 
b[40359] == 40359 && 
b[40360] == 40360 && 
b[40361] == 40361 && 
b[40362] == 40362 && 
b[40363] == 40363 && 
b[40364] == 40364 && 
b[40365] == 40365 && 
b[40366] == 40366 && 
b[40367] == 40367 && 
b[40368] == 40368 && 
b[40369] == 40369 && 
b[40370] == 40370 && 
b[40371] == 40371 && 
b[40372] == 40372 && 
b[40373] == 40373 && 
b[40374] == 40374 && 
b[40375] == 40375 && 
b[40376] == 40376 && 
b[40377] == 40377 && 
b[40378] == 40378 && 
b[40379] == 40379 && 
b[40380] == 40380 && 
b[40381] == 40381 && 
b[40382] == 40382 && 
b[40383] == 40383 && 
b[40384] == 40384 && 
b[40385] == 40385 && 
b[40386] == 40386 && 
b[40387] == 40387 && 
b[40388] == 40388 && 
b[40389] == 40389 && 
b[40390] == 40390 && 
b[40391] == 40391 && 
b[40392] == 40392 && 
b[40393] == 40393 && 
b[40394] == 40394 && 
b[40395] == 40395 && 
b[40396] == 40396 && 
b[40397] == 40397 && 
b[40398] == 40398 && 
b[40399] == 40399 && 
b[40400] == 40400 && 
b[40401] == 40401 && 
b[40402] == 40402 && 
b[40403] == 40403 && 
b[40404] == 40404 && 
b[40405] == 40405 && 
b[40406] == 40406 && 
b[40407] == 40407 && 
b[40408] == 40408 && 
b[40409] == 40409 && 
b[40410] == 40410 && 
b[40411] == 40411 && 
b[40412] == 40412 && 
b[40413] == 40413 && 
b[40414] == 40414 && 
b[40415] == 40415 && 
b[40416] == 40416 && 
b[40417] == 40417 && 
b[40418] == 40418 && 
b[40419] == 40419 && 
b[40420] == 40420 && 
b[40421] == 40421 && 
b[40422] == 40422 && 
b[40423] == 40423 && 
b[40424] == 40424 && 
b[40425] == 40425 && 
b[40426] == 40426 && 
b[40427] == 40427 && 
b[40428] == 40428 && 
b[40429] == 40429 && 
b[40430] == 40430 && 
b[40431] == 40431 && 
b[40432] == 40432 && 
b[40433] == 40433 && 
b[40434] == 40434 && 
b[40435] == 40435 && 
b[40436] == 40436 && 
b[40437] == 40437 && 
b[40438] == 40438 && 
b[40439] == 40439 && 
b[40440] == 40440 && 
b[40441] == 40441 && 
b[40442] == 40442 && 
b[40443] == 40443 && 
b[40444] == 40444 && 
b[40445] == 40445 && 
b[40446] == 40446 && 
b[40447] == 40447 && 
b[40448] == 40448 && 
b[40449] == 40449 && 
b[40450] == 40450 && 
b[40451] == 40451 && 
b[40452] == 40452 && 
b[40453] == 40453 && 
b[40454] == 40454 && 
b[40455] == 40455 && 
b[40456] == 40456 && 
b[40457] == 40457 && 
b[40458] == 40458 && 
b[40459] == 40459 && 
b[40460] == 40460 && 
b[40461] == 40461 && 
b[40462] == 40462 && 
b[40463] == 40463 && 
b[40464] == 40464 && 
b[40465] == 40465 && 
b[40466] == 40466 && 
b[40467] == 40467 && 
b[40468] == 40468 && 
b[40469] == 40469 && 
b[40470] == 40470 && 
b[40471] == 40471 && 
b[40472] == 40472 && 
b[40473] == 40473 && 
b[40474] == 40474 && 
b[40475] == 40475 && 
b[40476] == 40476 && 
b[40477] == 40477 && 
b[40478] == 40478 && 
b[40479] == 40479 && 
b[40480] == 40480 && 
b[40481] == 40481 && 
b[40482] == 40482 && 
b[40483] == 40483 && 
b[40484] == 40484 && 
b[40485] == 40485 && 
b[40486] == 40486 && 
b[40487] == 40487 && 
b[40488] == 40488 && 
b[40489] == 40489 && 
b[40490] == 40490 && 
b[40491] == 40491 && 
b[40492] == 40492 && 
b[40493] == 40493 && 
b[40494] == 40494 && 
b[40495] == 40495 && 
b[40496] == 40496 && 
b[40497] == 40497 && 
b[40498] == 40498 && 
b[40499] == 40499 && 
b[40500] == 40500 && 
b[40501] == 40501 && 
b[40502] == 40502 && 
b[40503] == 40503 && 
b[40504] == 40504 && 
b[40505] == 40505 && 
b[40506] == 40506 && 
b[40507] == 40507 && 
b[40508] == 40508 && 
b[40509] == 40509 && 
b[40510] == 40510 && 
b[40511] == 40511 && 
b[40512] == 40512 && 
b[40513] == 40513 && 
b[40514] == 40514 && 
b[40515] == 40515 && 
b[40516] == 40516 && 
b[40517] == 40517 && 
b[40518] == 40518 && 
b[40519] == 40519 && 
b[40520] == 40520 && 
b[40521] == 40521 && 
b[40522] == 40522 && 
b[40523] == 40523 && 
b[40524] == 40524 && 
b[40525] == 40525 && 
b[40526] == 40526 && 
b[40527] == 40527 && 
b[40528] == 40528 && 
b[40529] == 40529 && 
b[40530] == 40530 && 
b[40531] == 40531 && 
b[40532] == 40532 && 
b[40533] == 40533 && 
b[40534] == 40534 && 
b[40535] == 40535 && 
b[40536] == 40536 && 
b[40537] == 40537 && 
b[40538] == 40538 && 
b[40539] == 40539 && 
b[40540] == 40540 && 
b[40541] == 40541 && 
b[40542] == 40542 && 
b[40543] == 40543 && 
b[40544] == 40544 && 
b[40545] == 40545 && 
b[40546] == 40546 && 
b[40547] == 40547 && 
b[40548] == 40548 && 
b[40549] == 40549 && 
b[40550] == 40550 && 
b[40551] == 40551 && 
b[40552] == 40552 && 
b[40553] == 40553 && 
b[40554] == 40554 && 
b[40555] == 40555 && 
b[40556] == 40556 && 
b[40557] == 40557 && 
b[40558] == 40558 && 
b[40559] == 40559 && 
b[40560] == 40560 && 
b[40561] == 40561 && 
b[40562] == 40562 && 
b[40563] == 40563 && 
b[40564] == 40564 && 
b[40565] == 40565 && 
b[40566] == 40566 && 
b[40567] == 40567 && 
b[40568] == 40568 && 
b[40569] == 40569 && 
b[40570] == 40570 && 
b[40571] == 40571 && 
b[40572] == 40572 && 
b[40573] == 40573 && 
b[40574] == 40574 && 
b[40575] == 40575 && 
b[40576] == 40576 && 
b[40577] == 40577 && 
b[40578] == 40578 && 
b[40579] == 40579 && 
b[40580] == 40580 && 
b[40581] == 40581 && 
b[40582] == 40582 && 
b[40583] == 40583 && 
b[40584] == 40584 && 
b[40585] == 40585 && 
b[40586] == 40586 && 
b[40587] == 40587 && 
b[40588] == 40588 && 
b[40589] == 40589 && 
b[40590] == 40590 && 
b[40591] == 40591 && 
b[40592] == 40592 && 
b[40593] == 40593 && 
b[40594] == 40594 && 
b[40595] == 40595 && 
b[40596] == 40596 && 
b[40597] == 40597 && 
b[40598] == 40598 && 
b[40599] == 40599 && 
b[40600] == 40600 && 
b[40601] == 40601 && 
b[40602] == 40602 && 
b[40603] == 40603 && 
b[40604] == 40604 && 
b[40605] == 40605 && 
b[40606] == 40606 && 
b[40607] == 40607 && 
b[40608] == 40608 && 
b[40609] == 40609 && 
b[40610] == 40610 && 
b[40611] == 40611 && 
b[40612] == 40612 && 
b[40613] == 40613 && 
b[40614] == 40614 && 
b[40615] == 40615 && 
b[40616] == 40616 && 
b[40617] == 40617 && 
b[40618] == 40618 && 
b[40619] == 40619 && 
b[40620] == 40620 && 
b[40621] == 40621 && 
b[40622] == 40622 && 
b[40623] == 40623 && 
b[40624] == 40624 && 
b[40625] == 40625 && 
b[40626] == 40626 && 
b[40627] == 40627 && 
b[40628] == 40628 && 
b[40629] == 40629 && 
b[40630] == 40630 && 
b[40631] == 40631 && 
b[40632] == 40632 && 
b[40633] == 40633 && 
b[40634] == 40634 && 
b[40635] == 40635 && 
b[40636] == 40636 && 
b[40637] == 40637 && 
b[40638] == 40638 && 
b[40639] == 40639 && 
b[40640] == 40640 && 
b[40641] == 40641 && 
b[40642] == 40642 && 
b[40643] == 40643 && 
b[40644] == 40644 && 
b[40645] == 40645 && 
b[40646] == 40646 && 
b[40647] == 40647 && 
b[40648] == 40648 && 
b[40649] == 40649 && 
b[40650] == 40650 && 
b[40651] == 40651 && 
b[40652] == 40652 && 
b[40653] == 40653 && 
b[40654] == 40654 && 
b[40655] == 40655 && 
b[40656] == 40656 && 
b[40657] == 40657 && 
b[40658] == 40658 && 
b[40659] == 40659 && 
b[40660] == 40660 && 
b[40661] == 40661 && 
b[40662] == 40662 && 
b[40663] == 40663 && 
b[40664] == 40664 && 
b[40665] == 40665 && 
b[40666] == 40666 && 
b[40667] == 40667 && 
b[40668] == 40668 && 
b[40669] == 40669 && 
b[40670] == 40670 && 
b[40671] == 40671 && 
b[40672] == 40672 && 
b[40673] == 40673 && 
b[40674] == 40674 && 
b[40675] == 40675 && 
b[40676] == 40676 && 
b[40677] == 40677 && 
b[40678] == 40678 && 
b[40679] == 40679 && 
b[40680] == 40680 && 
b[40681] == 40681 && 
b[40682] == 40682 && 
b[40683] == 40683 && 
b[40684] == 40684 && 
b[40685] == 40685 && 
b[40686] == 40686 && 
b[40687] == 40687 && 
b[40688] == 40688 && 
b[40689] == 40689 && 
b[40690] == 40690 && 
b[40691] == 40691 && 
b[40692] == 40692 && 
b[40693] == 40693 && 
b[40694] == 40694 && 
b[40695] == 40695 && 
b[40696] == 40696 && 
b[40697] == 40697 && 
b[40698] == 40698 && 
b[40699] == 40699 && 
b[40700] == 40700 && 
b[40701] == 40701 && 
b[40702] == 40702 && 
b[40703] == 40703 && 
b[40704] == 40704 && 
b[40705] == 40705 && 
b[40706] == 40706 && 
b[40707] == 40707 && 
b[40708] == 40708 && 
b[40709] == 40709 && 
b[40710] == 40710 && 
b[40711] == 40711 && 
b[40712] == 40712 && 
b[40713] == 40713 && 
b[40714] == 40714 && 
b[40715] == 40715 && 
b[40716] == 40716 && 
b[40717] == 40717 && 
b[40718] == 40718 && 
b[40719] == 40719 && 
b[40720] == 40720 && 
b[40721] == 40721 && 
b[40722] == 40722 && 
b[40723] == 40723 && 
b[40724] == 40724 && 
b[40725] == 40725 && 
b[40726] == 40726 && 
b[40727] == 40727 && 
b[40728] == 40728 && 
b[40729] == 40729 && 
b[40730] == 40730 && 
b[40731] == 40731 && 
b[40732] == 40732 && 
b[40733] == 40733 && 
b[40734] == 40734 && 
b[40735] == 40735 && 
b[40736] == 40736 && 
b[40737] == 40737 && 
b[40738] == 40738 && 
b[40739] == 40739 && 
b[40740] == 40740 && 
b[40741] == 40741 && 
b[40742] == 40742 && 
b[40743] == 40743 && 
b[40744] == 40744 && 
b[40745] == 40745 && 
b[40746] == 40746 && 
b[40747] == 40747 && 
b[40748] == 40748 && 
b[40749] == 40749 && 
b[40750] == 40750 && 
b[40751] == 40751 && 
b[40752] == 40752 && 
b[40753] == 40753 && 
b[40754] == 40754 && 
b[40755] == 40755 && 
b[40756] == 40756 && 
b[40757] == 40757 && 
b[40758] == 40758 && 
b[40759] == 40759 && 
b[40760] == 40760 && 
b[40761] == 40761 && 
b[40762] == 40762 && 
b[40763] == 40763 && 
b[40764] == 40764 && 
b[40765] == 40765 && 
b[40766] == 40766 && 
b[40767] == 40767 && 
b[40768] == 40768 && 
b[40769] == 40769 && 
b[40770] == 40770 && 
b[40771] == 40771 && 
b[40772] == 40772 && 
b[40773] == 40773 && 
b[40774] == 40774 && 
b[40775] == 40775 && 
b[40776] == 40776 && 
b[40777] == 40777 && 
b[40778] == 40778 && 
b[40779] == 40779 && 
b[40780] == 40780 && 
b[40781] == 40781 && 
b[40782] == 40782 && 
b[40783] == 40783 && 
b[40784] == 40784 && 
b[40785] == 40785 && 
b[40786] == 40786 && 
b[40787] == 40787 && 
b[40788] == 40788 && 
b[40789] == 40789 && 
b[40790] == 40790 && 
b[40791] == 40791 && 
b[40792] == 40792 && 
b[40793] == 40793 && 
b[40794] == 40794 && 
b[40795] == 40795 && 
b[40796] == 40796 && 
b[40797] == 40797 && 
b[40798] == 40798 && 
b[40799] == 40799 && 
b[40800] == 40800 && 
b[40801] == 40801 && 
b[40802] == 40802 && 
b[40803] == 40803 && 
b[40804] == 40804 && 
b[40805] == 40805 && 
b[40806] == 40806 && 
b[40807] == 40807 && 
b[40808] == 40808 && 
b[40809] == 40809 && 
b[40810] == 40810 && 
b[40811] == 40811 && 
b[40812] == 40812 && 
b[40813] == 40813 && 
b[40814] == 40814 && 
b[40815] == 40815 && 
b[40816] == 40816 && 
b[40817] == 40817 && 
b[40818] == 40818 && 
b[40819] == 40819 && 
b[40820] == 40820 && 
b[40821] == 40821 && 
b[40822] == 40822 && 
b[40823] == 40823 && 
b[40824] == 40824 && 
b[40825] == 40825 && 
b[40826] == 40826 && 
b[40827] == 40827 && 
b[40828] == 40828 && 
b[40829] == 40829 && 
b[40830] == 40830 && 
b[40831] == 40831 && 
b[40832] == 40832 && 
b[40833] == 40833 && 
b[40834] == 40834 && 
b[40835] == 40835 && 
b[40836] == 40836 && 
b[40837] == 40837 && 
b[40838] == 40838 && 
b[40839] == 40839 && 
b[40840] == 40840 && 
b[40841] == 40841 && 
b[40842] == 40842 && 
b[40843] == 40843 && 
b[40844] == 40844 && 
b[40845] == 40845 && 
b[40846] == 40846 && 
b[40847] == 40847 && 
b[40848] == 40848 && 
b[40849] == 40849 && 
b[40850] == 40850 && 
b[40851] == 40851 && 
b[40852] == 40852 && 
b[40853] == 40853 && 
b[40854] == 40854 && 
b[40855] == 40855 && 
b[40856] == 40856 && 
b[40857] == 40857 && 
b[40858] == 40858 && 
b[40859] == 40859 && 
b[40860] == 40860 && 
b[40861] == 40861 && 
b[40862] == 40862 && 
b[40863] == 40863 && 
b[40864] == 40864 && 
b[40865] == 40865 && 
b[40866] == 40866 && 
b[40867] == 40867 && 
b[40868] == 40868 && 
b[40869] == 40869 && 
b[40870] == 40870 && 
b[40871] == 40871 && 
b[40872] == 40872 && 
b[40873] == 40873 && 
b[40874] == 40874 && 
b[40875] == 40875 && 
b[40876] == 40876 && 
b[40877] == 40877 && 
b[40878] == 40878 && 
b[40879] == 40879 && 
b[40880] == 40880 && 
b[40881] == 40881 && 
b[40882] == 40882 && 
b[40883] == 40883 && 
b[40884] == 40884 && 
b[40885] == 40885 && 
b[40886] == 40886 && 
b[40887] == 40887 && 
b[40888] == 40888 && 
b[40889] == 40889 && 
b[40890] == 40890 && 
b[40891] == 40891 && 
b[40892] == 40892 && 
b[40893] == 40893 && 
b[40894] == 40894 && 
b[40895] == 40895 && 
b[40896] == 40896 && 
b[40897] == 40897 && 
b[40898] == 40898 && 
b[40899] == 40899 && 
b[40900] == 40900 && 
b[40901] == 40901 && 
b[40902] == 40902 && 
b[40903] == 40903 && 
b[40904] == 40904 && 
b[40905] == 40905 && 
b[40906] == 40906 && 
b[40907] == 40907 && 
b[40908] == 40908 && 
b[40909] == 40909 && 
b[40910] == 40910 && 
b[40911] == 40911 && 
b[40912] == 40912 && 
b[40913] == 40913 && 
b[40914] == 40914 && 
b[40915] == 40915 && 
b[40916] == 40916 && 
b[40917] == 40917 && 
b[40918] == 40918 && 
b[40919] == 40919 && 
b[40920] == 40920 && 
b[40921] == 40921 && 
b[40922] == 40922 && 
b[40923] == 40923 && 
b[40924] == 40924 && 
b[40925] == 40925 && 
b[40926] == 40926 && 
b[40927] == 40927 && 
b[40928] == 40928 && 
b[40929] == 40929 && 
b[40930] == 40930 && 
b[40931] == 40931 && 
b[40932] == 40932 && 
b[40933] == 40933 && 
b[40934] == 40934 && 
b[40935] == 40935 && 
b[40936] == 40936 && 
b[40937] == 40937 && 
b[40938] == 40938 && 
b[40939] == 40939 && 
b[40940] == 40940 && 
b[40941] == 40941 && 
b[40942] == 40942 && 
b[40943] == 40943 && 
b[40944] == 40944 && 
b[40945] == 40945 && 
b[40946] == 40946 && 
b[40947] == 40947 && 
b[40948] == 40948 && 
b[40949] == 40949 && 
b[40950] == 40950 && 
b[40951] == 40951 && 
b[40952] == 40952 && 
b[40953] == 40953 && 
b[40954] == 40954 && 
b[40955] == 40955 && 
b[40956] == 40956 && 
b[40957] == 40957 && 
b[40958] == 40958 && 
b[40959] == 40959 && 
b[40960] == 40960 && 
b[40961] == 40961 && 
b[40962] == 40962 && 
b[40963] == 40963 && 
b[40964] == 40964 && 
b[40965] == 40965 && 
b[40966] == 40966 && 
b[40967] == 40967 && 
b[40968] == 40968 && 
b[40969] == 40969 && 
b[40970] == 40970 && 
b[40971] == 40971 && 
b[40972] == 40972 && 
b[40973] == 40973 && 
b[40974] == 40974 && 
b[40975] == 40975 && 
b[40976] == 40976 && 
b[40977] == 40977 && 
b[40978] == 40978 && 
b[40979] == 40979 && 
b[40980] == 40980 && 
b[40981] == 40981 && 
b[40982] == 40982 && 
b[40983] == 40983 && 
b[40984] == 40984 && 
b[40985] == 40985 && 
b[40986] == 40986 && 
b[40987] == 40987 && 
b[40988] == 40988 && 
b[40989] == 40989 && 
b[40990] == 40990 && 
b[40991] == 40991 && 
b[40992] == 40992 && 
b[40993] == 40993 && 
b[40994] == 40994 && 
b[40995] == 40995 && 
b[40996] == 40996 && 
b[40997] == 40997 && 
b[40998] == 40998 && 
b[40999] == 40999 && 
b[41000] == 41000 && 
b[41001] == 41001 && 
b[41002] == 41002 && 
b[41003] == 41003 && 
b[41004] == 41004 && 
b[41005] == 41005 && 
b[41006] == 41006 && 
b[41007] == 41007 && 
b[41008] == 41008 && 
b[41009] == 41009 && 
b[41010] == 41010 && 
b[41011] == 41011 && 
b[41012] == 41012 && 
b[41013] == 41013 && 
b[41014] == 41014 && 
b[41015] == 41015 && 
b[41016] == 41016 && 
b[41017] == 41017 && 
b[41018] == 41018 && 
b[41019] == 41019 && 
b[41020] == 41020 && 
b[41021] == 41021 && 
b[41022] == 41022 && 
b[41023] == 41023 && 
b[41024] == 41024 && 
b[41025] == 41025 && 
b[41026] == 41026 && 
b[41027] == 41027 && 
b[41028] == 41028 && 
b[41029] == 41029 && 
b[41030] == 41030 && 
b[41031] == 41031 && 
b[41032] == 41032 && 
b[41033] == 41033 && 
b[41034] == 41034 && 
b[41035] == 41035 && 
b[41036] == 41036 && 
b[41037] == 41037 && 
b[41038] == 41038 && 
b[41039] == 41039 && 
b[41040] == 41040 && 
b[41041] == 41041 && 
b[41042] == 41042 && 
b[41043] == 41043 && 
b[41044] == 41044 && 
b[41045] == 41045 && 
b[41046] == 41046 && 
b[41047] == 41047 && 
b[41048] == 41048 && 
b[41049] == 41049 && 
b[41050] == 41050 && 
b[41051] == 41051 && 
b[41052] == 41052 && 
b[41053] == 41053 && 
b[41054] == 41054 && 
b[41055] == 41055 && 
b[41056] == 41056 && 
b[41057] == 41057 && 
b[41058] == 41058 && 
b[41059] == 41059 && 
b[41060] == 41060 && 
b[41061] == 41061 && 
b[41062] == 41062 && 
b[41063] == 41063 && 
b[41064] == 41064 && 
b[41065] == 41065 && 
b[41066] == 41066 && 
b[41067] == 41067 && 
b[41068] == 41068 && 
b[41069] == 41069 && 
b[41070] == 41070 && 
b[41071] == 41071 && 
b[41072] == 41072 && 
b[41073] == 41073 && 
b[41074] == 41074 && 
b[41075] == 41075 && 
b[41076] == 41076 && 
b[41077] == 41077 && 
b[41078] == 41078 && 
b[41079] == 41079 && 
b[41080] == 41080 && 
b[41081] == 41081 && 
b[41082] == 41082 && 
b[41083] == 41083 && 
b[41084] == 41084 && 
b[41085] == 41085 && 
b[41086] == 41086 && 
b[41087] == 41087 && 
b[41088] == 41088 && 
b[41089] == 41089 && 
b[41090] == 41090 && 
b[41091] == 41091 && 
b[41092] == 41092 && 
b[41093] == 41093 && 
b[41094] == 41094 && 
b[41095] == 41095 && 
b[41096] == 41096 && 
b[41097] == 41097 && 
b[41098] == 41098 && 
b[41099] == 41099 && 
b[41100] == 41100 && 
b[41101] == 41101 && 
b[41102] == 41102 && 
b[41103] == 41103 && 
b[41104] == 41104 && 
b[41105] == 41105 && 
b[41106] == 41106 && 
b[41107] == 41107 && 
b[41108] == 41108 && 
b[41109] == 41109 && 
b[41110] == 41110 && 
b[41111] == 41111 && 
b[41112] == 41112 && 
b[41113] == 41113 && 
b[41114] == 41114 && 
b[41115] == 41115 && 
b[41116] == 41116 && 
b[41117] == 41117 && 
b[41118] == 41118 && 
b[41119] == 41119 && 
b[41120] == 41120 && 
b[41121] == 41121 && 
b[41122] == 41122 && 
b[41123] == 41123 && 
b[41124] == 41124 && 
b[41125] == 41125 && 
b[41126] == 41126 && 
b[41127] == 41127 && 
b[41128] == 41128 && 
b[41129] == 41129 && 
b[41130] == 41130 && 
b[41131] == 41131 && 
b[41132] == 41132 && 
b[41133] == 41133 && 
b[41134] == 41134 && 
b[41135] == 41135 && 
b[41136] == 41136 && 
b[41137] == 41137 && 
b[41138] == 41138 && 
b[41139] == 41139 && 
b[41140] == 41140 && 
b[41141] == 41141 && 
b[41142] == 41142 && 
b[41143] == 41143 && 
b[41144] == 41144 && 
b[41145] == 41145 && 
b[41146] == 41146 && 
b[41147] == 41147 && 
b[41148] == 41148 && 
b[41149] == 41149 && 
b[41150] == 41150 && 
b[41151] == 41151 && 
b[41152] == 41152 && 
b[41153] == 41153 && 
b[41154] == 41154 && 
b[41155] == 41155 && 
b[41156] == 41156 && 
b[41157] == 41157 && 
b[41158] == 41158 && 
b[41159] == 41159 && 
b[41160] == 41160 && 
b[41161] == 41161 && 
b[41162] == 41162 && 
b[41163] == 41163 && 
b[41164] == 41164 && 
b[41165] == 41165 && 
b[41166] == 41166 && 
b[41167] == 41167 && 
b[41168] == 41168 && 
b[41169] == 41169 && 
b[41170] == 41170 && 
b[41171] == 41171 && 
b[41172] == 41172 && 
b[41173] == 41173 && 
b[41174] == 41174 && 
b[41175] == 41175 && 
b[41176] == 41176 && 
b[41177] == 41177 && 
b[41178] == 41178 && 
b[41179] == 41179 && 
b[41180] == 41180 && 
b[41181] == 41181 && 
b[41182] == 41182 && 
b[41183] == 41183 && 
b[41184] == 41184 && 
b[41185] == 41185 && 
b[41186] == 41186 && 
b[41187] == 41187 && 
b[41188] == 41188 && 
b[41189] == 41189 && 
b[41190] == 41190 && 
b[41191] == 41191 && 
b[41192] == 41192 && 
b[41193] == 41193 && 
b[41194] == 41194 && 
b[41195] == 41195 && 
b[41196] == 41196 && 
b[41197] == 41197 && 
b[41198] == 41198 && 
b[41199] == 41199 && 
b[41200] == 41200 && 
b[41201] == 41201 && 
b[41202] == 41202 && 
b[41203] == 41203 && 
b[41204] == 41204 && 
b[41205] == 41205 && 
b[41206] == 41206 && 
b[41207] == 41207 && 
b[41208] == 41208 && 
b[41209] == 41209 && 
b[41210] == 41210 && 
b[41211] == 41211 && 
b[41212] == 41212 && 
b[41213] == 41213 && 
b[41214] == 41214 && 
b[41215] == 41215 && 
b[41216] == 41216 && 
b[41217] == 41217 && 
b[41218] == 41218 && 
b[41219] == 41219 && 
b[41220] == 41220 && 
b[41221] == 41221 && 
b[41222] == 41222 && 
b[41223] == 41223 && 
b[41224] == 41224 && 
b[41225] == 41225 && 
b[41226] == 41226 && 
b[41227] == 41227 && 
b[41228] == 41228 && 
b[41229] == 41229 && 
b[41230] == 41230 && 
b[41231] == 41231 && 
b[41232] == 41232 && 
b[41233] == 41233 && 
b[41234] == 41234 && 
b[41235] == 41235 && 
b[41236] == 41236 && 
b[41237] == 41237 && 
b[41238] == 41238 && 
b[41239] == 41239 && 
b[41240] == 41240 && 
b[41241] == 41241 && 
b[41242] == 41242 && 
b[41243] == 41243 && 
b[41244] == 41244 && 
b[41245] == 41245 && 
b[41246] == 41246 && 
b[41247] == 41247 && 
b[41248] == 41248 && 
b[41249] == 41249 && 
b[41250] == 41250 && 
b[41251] == 41251 && 
b[41252] == 41252 && 
b[41253] == 41253 && 
b[41254] == 41254 && 
b[41255] == 41255 && 
b[41256] == 41256 && 
b[41257] == 41257 && 
b[41258] == 41258 && 
b[41259] == 41259 && 
b[41260] == 41260 && 
b[41261] == 41261 && 
b[41262] == 41262 && 
b[41263] == 41263 && 
b[41264] == 41264 && 
b[41265] == 41265 && 
b[41266] == 41266 && 
b[41267] == 41267 && 
b[41268] == 41268 && 
b[41269] == 41269 && 
b[41270] == 41270 && 
b[41271] == 41271 && 
b[41272] == 41272 && 
b[41273] == 41273 && 
b[41274] == 41274 && 
b[41275] == 41275 && 
b[41276] == 41276 && 
b[41277] == 41277 && 
b[41278] == 41278 && 
b[41279] == 41279 && 
b[41280] == 41280 && 
b[41281] == 41281 && 
b[41282] == 41282 && 
b[41283] == 41283 && 
b[41284] == 41284 && 
b[41285] == 41285 && 
b[41286] == 41286 && 
b[41287] == 41287 && 
b[41288] == 41288 && 
b[41289] == 41289 && 
b[41290] == 41290 && 
b[41291] == 41291 && 
b[41292] == 41292 && 
b[41293] == 41293 && 
b[41294] == 41294 && 
b[41295] == 41295 && 
b[41296] == 41296 && 
b[41297] == 41297 && 
b[41298] == 41298 && 
b[41299] == 41299 && 
b[41300] == 41300 && 
b[41301] == 41301 && 
b[41302] == 41302 && 
b[41303] == 41303 && 
b[41304] == 41304 && 
b[41305] == 41305 && 
b[41306] == 41306 && 
b[41307] == 41307 && 
b[41308] == 41308 && 
b[41309] == 41309 && 
b[41310] == 41310 && 
b[41311] == 41311 && 
b[41312] == 41312 && 
b[41313] == 41313 && 
b[41314] == 41314 && 
b[41315] == 41315 && 
b[41316] == 41316 && 
b[41317] == 41317 && 
b[41318] == 41318 && 
b[41319] == 41319 && 
b[41320] == 41320 && 
b[41321] == 41321 && 
b[41322] == 41322 && 
b[41323] == 41323 && 
b[41324] == 41324 && 
b[41325] == 41325 && 
b[41326] == 41326 && 
b[41327] == 41327 && 
b[41328] == 41328 && 
b[41329] == 41329 && 
b[41330] == 41330 && 
b[41331] == 41331 && 
b[41332] == 41332 && 
b[41333] == 41333 && 
b[41334] == 41334 && 
b[41335] == 41335 && 
b[41336] == 41336 && 
b[41337] == 41337 && 
b[41338] == 41338 && 
b[41339] == 41339 && 
b[41340] == 41340 && 
b[41341] == 41341 && 
b[41342] == 41342 && 
b[41343] == 41343 && 
b[41344] == 41344 && 
b[41345] == 41345 && 
b[41346] == 41346 && 
b[41347] == 41347 && 
b[41348] == 41348 && 
b[41349] == 41349 && 
b[41350] == 41350 && 
b[41351] == 41351 && 
b[41352] == 41352 && 
b[41353] == 41353 && 
b[41354] == 41354 && 
b[41355] == 41355 && 
b[41356] == 41356 && 
b[41357] == 41357 && 
b[41358] == 41358 && 
b[41359] == 41359 && 
b[41360] == 41360 && 
b[41361] == 41361 && 
b[41362] == 41362 && 
b[41363] == 41363 && 
b[41364] == 41364 && 
b[41365] == 41365 && 
b[41366] == 41366 && 
b[41367] == 41367 && 
b[41368] == 41368 && 
b[41369] == 41369 && 
b[41370] == 41370 && 
b[41371] == 41371 && 
b[41372] == 41372 && 
b[41373] == 41373 && 
b[41374] == 41374 && 
b[41375] == 41375 && 
b[41376] == 41376 && 
b[41377] == 41377 && 
b[41378] == 41378 && 
b[41379] == 41379 && 
b[41380] == 41380 && 
b[41381] == 41381 && 
b[41382] == 41382 && 
b[41383] == 41383 && 
b[41384] == 41384 && 
b[41385] == 41385 && 
b[41386] == 41386 && 
b[41387] == 41387 && 
b[41388] == 41388 && 
b[41389] == 41389 && 
b[41390] == 41390 && 
b[41391] == 41391 && 
b[41392] == 41392 && 
b[41393] == 41393 && 
b[41394] == 41394 && 
b[41395] == 41395 && 
b[41396] == 41396 && 
b[41397] == 41397 && 
b[41398] == 41398 && 
b[41399] == 41399 && 
b[41400] == 41400 && 
b[41401] == 41401 && 
b[41402] == 41402 && 
b[41403] == 41403 && 
b[41404] == 41404 && 
b[41405] == 41405 && 
b[41406] == 41406 && 
b[41407] == 41407 && 
b[41408] == 41408 && 
b[41409] == 41409 && 
b[41410] == 41410 && 
b[41411] == 41411 && 
b[41412] == 41412 && 
b[41413] == 41413 && 
b[41414] == 41414 && 
b[41415] == 41415 && 
b[41416] == 41416 && 
b[41417] == 41417 && 
b[41418] == 41418 && 
b[41419] == 41419 && 
b[41420] == 41420 && 
b[41421] == 41421 && 
b[41422] == 41422 && 
b[41423] == 41423 && 
b[41424] == 41424 && 
b[41425] == 41425 && 
b[41426] == 41426 && 
b[41427] == 41427 && 
b[41428] == 41428 && 
b[41429] == 41429 && 
b[41430] == 41430 && 
b[41431] == 41431 && 
b[41432] == 41432 && 
b[41433] == 41433 && 
b[41434] == 41434 && 
b[41435] == 41435 && 
b[41436] == 41436 && 
b[41437] == 41437 && 
b[41438] == 41438 && 
b[41439] == 41439 && 
b[41440] == 41440 && 
b[41441] == 41441 && 
b[41442] == 41442 && 
b[41443] == 41443 && 
b[41444] == 41444 && 
b[41445] == 41445 && 
b[41446] == 41446 && 
b[41447] == 41447 && 
b[41448] == 41448 && 
b[41449] == 41449 && 
b[41450] == 41450 && 
b[41451] == 41451 && 
b[41452] == 41452 && 
b[41453] == 41453 && 
b[41454] == 41454 && 
b[41455] == 41455 && 
b[41456] == 41456 && 
b[41457] == 41457 && 
b[41458] == 41458 && 
b[41459] == 41459 && 
b[41460] == 41460 && 
b[41461] == 41461 && 
b[41462] == 41462 && 
b[41463] == 41463 && 
b[41464] == 41464 && 
b[41465] == 41465 && 
b[41466] == 41466 && 
b[41467] == 41467 && 
b[41468] == 41468 && 
b[41469] == 41469 && 
b[41470] == 41470 && 
b[41471] == 41471 && 
b[41472] == 41472 && 
b[41473] == 41473 && 
b[41474] == 41474 && 
b[41475] == 41475 && 
b[41476] == 41476 && 
b[41477] == 41477 && 
b[41478] == 41478 && 
b[41479] == 41479 && 
b[41480] == 41480 && 
b[41481] == 41481 && 
b[41482] == 41482 && 
b[41483] == 41483 && 
b[41484] == 41484 && 
b[41485] == 41485 && 
b[41486] == 41486 && 
b[41487] == 41487 && 
b[41488] == 41488 && 
b[41489] == 41489 && 
b[41490] == 41490 && 
b[41491] == 41491 && 
b[41492] == 41492 && 
b[41493] == 41493 && 
b[41494] == 41494 && 
b[41495] == 41495 && 
b[41496] == 41496 && 
b[41497] == 41497 && 
b[41498] == 41498 && 
b[41499] == 41499 && 
b[41500] == 41500 && 
b[41501] == 41501 && 
b[41502] == 41502 && 
b[41503] == 41503 && 
b[41504] == 41504 && 
b[41505] == 41505 && 
b[41506] == 41506 && 
b[41507] == 41507 && 
b[41508] == 41508 && 
b[41509] == 41509 && 
b[41510] == 41510 && 
b[41511] == 41511 && 
b[41512] == 41512 && 
b[41513] == 41513 && 
b[41514] == 41514 && 
b[41515] == 41515 && 
b[41516] == 41516 && 
b[41517] == 41517 && 
b[41518] == 41518 && 
b[41519] == 41519 && 
b[41520] == 41520 && 
b[41521] == 41521 && 
b[41522] == 41522 && 
b[41523] == 41523 && 
b[41524] == 41524 && 
b[41525] == 41525 && 
b[41526] == 41526 && 
b[41527] == 41527 && 
b[41528] == 41528 && 
b[41529] == 41529 && 
b[41530] == 41530 && 
b[41531] == 41531 && 
b[41532] == 41532 && 
b[41533] == 41533 && 
b[41534] == 41534 && 
b[41535] == 41535 && 
b[41536] == 41536 && 
b[41537] == 41537 && 
b[41538] == 41538 && 
b[41539] == 41539 && 
b[41540] == 41540 && 
b[41541] == 41541 && 
b[41542] == 41542 && 
b[41543] == 41543 && 
b[41544] == 41544 && 
b[41545] == 41545 && 
b[41546] == 41546 && 
b[41547] == 41547 && 
b[41548] == 41548 && 
b[41549] == 41549 && 
b[41550] == 41550 && 
b[41551] == 41551 && 
b[41552] == 41552 && 
b[41553] == 41553 && 
b[41554] == 41554 && 
b[41555] == 41555 && 
b[41556] == 41556 && 
b[41557] == 41557 && 
b[41558] == 41558 && 
b[41559] == 41559 && 
b[41560] == 41560 && 
b[41561] == 41561 && 
b[41562] == 41562 && 
b[41563] == 41563 && 
b[41564] == 41564 && 
b[41565] == 41565 && 
b[41566] == 41566 && 
b[41567] == 41567 && 
b[41568] == 41568 && 
b[41569] == 41569 && 
b[41570] == 41570 && 
b[41571] == 41571 && 
b[41572] == 41572 && 
b[41573] == 41573 && 
b[41574] == 41574 && 
b[41575] == 41575 && 
b[41576] == 41576 && 
b[41577] == 41577 && 
b[41578] == 41578 && 
b[41579] == 41579 && 
b[41580] == 41580 && 
b[41581] == 41581 && 
b[41582] == 41582 && 
b[41583] == 41583 && 
b[41584] == 41584 && 
b[41585] == 41585 && 
b[41586] == 41586 && 
b[41587] == 41587 && 
b[41588] == 41588 && 
b[41589] == 41589 && 
b[41590] == 41590 && 
b[41591] == 41591 && 
b[41592] == 41592 && 
b[41593] == 41593 && 
b[41594] == 41594 && 
b[41595] == 41595 && 
b[41596] == 41596 && 
b[41597] == 41597 && 
b[41598] == 41598 && 
b[41599] == 41599 && 
b[41600] == 41600 && 
b[41601] == 41601 && 
b[41602] == 41602 && 
b[41603] == 41603 && 
b[41604] == 41604 && 
b[41605] == 41605 && 
b[41606] == 41606 && 
b[41607] == 41607 && 
b[41608] == 41608 && 
b[41609] == 41609 && 
b[41610] == 41610 && 
b[41611] == 41611 && 
b[41612] == 41612 && 
b[41613] == 41613 && 
b[41614] == 41614 && 
b[41615] == 41615 && 
b[41616] == 41616 && 
b[41617] == 41617 && 
b[41618] == 41618 && 
b[41619] == 41619 && 
b[41620] == 41620 && 
b[41621] == 41621 && 
b[41622] == 41622 && 
b[41623] == 41623 && 
b[41624] == 41624 && 
b[41625] == 41625 && 
b[41626] == 41626 && 
b[41627] == 41627 && 
b[41628] == 41628 && 
b[41629] == 41629 && 
b[41630] == 41630 && 
b[41631] == 41631 && 
b[41632] == 41632 && 
b[41633] == 41633 && 
b[41634] == 41634 && 
b[41635] == 41635 && 
b[41636] == 41636 && 
b[41637] == 41637 && 
b[41638] == 41638 && 
b[41639] == 41639 && 
b[41640] == 41640 && 
b[41641] == 41641 && 
b[41642] == 41642 && 
b[41643] == 41643 && 
b[41644] == 41644 && 
b[41645] == 41645 && 
b[41646] == 41646 && 
b[41647] == 41647 && 
b[41648] == 41648 && 
b[41649] == 41649 && 
b[41650] == 41650 && 
b[41651] == 41651 && 
b[41652] == 41652 && 
b[41653] == 41653 && 
b[41654] == 41654 && 
b[41655] == 41655 && 
b[41656] == 41656 && 
b[41657] == 41657 && 
b[41658] == 41658 && 
b[41659] == 41659 && 
b[41660] == 41660 && 
b[41661] == 41661 && 
b[41662] == 41662 && 
b[41663] == 41663 && 
b[41664] == 41664 && 
b[41665] == 41665 && 
b[41666] == 41666 && 
b[41667] == 41667 && 
b[41668] == 41668 && 
b[41669] == 41669 && 
b[41670] == 41670 && 
b[41671] == 41671 && 
b[41672] == 41672 && 
b[41673] == 41673 && 
b[41674] == 41674 && 
b[41675] == 41675 && 
b[41676] == 41676 && 
b[41677] == 41677 && 
b[41678] == 41678 && 
b[41679] == 41679 && 
b[41680] == 41680 && 
b[41681] == 41681 && 
b[41682] == 41682 && 
b[41683] == 41683 && 
b[41684] == 41684 && 
b[41685] == 41685 && 
b[41686] == 41686 && 
b[41687] == 41687 && 
b[41688] == 41688 && 
b[41689] == 41689 && 
b[41690] == 41690 && 
b[41691] == 41691 && 
b[41692] == 41692 && 
b[41693] == 41693 && 
b[41694] == 41694 && 
b[41695] == 41695 && 
b[41696] == 41696 && 
b[41697] == 41697 && 
b[41698] == 41698 && 
b[41699] == 41699 && 
b[41700] == 41700 && 
b[41701] == 41701 && 
b[41702] == 41702 && 
b[41703] == 41703 && 
b[41704] == 41704 && 
b[41705] == 41705 && 
b[41706] == 41706 && 
b[41707] == 41707 && 
b[41708] == 41708 && 
b[41709] == 41709 && 
b[41710] == 41710 && 
b[41711] == 41711 && 
b[41712] == 41712 && 
b[41713] == 41713 && 
b[41714] == 41714 && 
b[41715] == 41715 && 
b[41716] == 41716 && 
b[41717] == 41717 && 
b[41718] == 41718 && 
b[41719] == 41719 && 
b[41720] == 41720 && 
b[41721] == 41721 && 
b[41722] == 41722 && 
b[41723] == 41723 && 
b[41724] == 41724 && 
b[41725] == 41725 && 
b[41726] == 41726 && 
b[41727] == 41727 && 
b[41728] == 41728 && 
b[41729] == 41729 && 
b[41730] == 41730 && 
b[41731] == 41731 && 
b[41732] == 41732 && 
b[41733] == 41733 && 
b[41734] == 41734 && 
b[41735] == 41735 && 
b[41736] == 41736 && 
b[41737] == 41737 && 
b[41738] == 41738 && 
b[41739] == 41739 && 
b[41740] == 41740 && 
b[41741] == 41741 && 
b[41742] == 41742 && 
b[41743] == 41743 && 
b[41744] == 41744 && 
b[41745] == 41745 && 
b[41746] == 41746 && 
b[41747] == 41747 && 
b[41748] == 41748 && 
b[41749] == 41749 && 
b[41750] == 41750 && 
b[41751] == 41751 && 
b[41752] == 41752 && 
b[41753] == 41753 && 
b[41754] == 41754 && 
b[41755] == 41755 && 
b[41756] == 41756 && 
b[41757] == 41757 && 
b[41758] == 41758 && 
b[41759] == 41759 && 
b[41760] == 41760 && 
b[41761] == 41761 && 
b[41762] == 41762 && 
b[41763] == 41763 && 
b[41764] == 41764 && 
b[41765] == 41765 && 
b[41766] == 41766 && 
b[41767] == 41767 && 
b[41768] == 41768 && 
b[41769] == 41769 && 
b[41770] == 41770 && 
b[41771] == 41771 && 
b[41772] == 41772 && 
b[41773] == 41773 && 
b[41774] == 41774 && 
b[41775] == 41775 && 
b[41776] == 41776 && 
b[41777] == 41777 && 
b[41778] == 41778 && 
b[41779] == 41779 && 
b[41780] == 41780 && 
b[41781] == 41781 && 
b[41782] == 41782 && 
b[41783] == 41783 && 
b[41784] == 41784 && 
b[41785] == 41785 && 
b[41786] == 41786 && 
b[41787] == 41787 && 
b[41788] == 41788 && 
b[41789] == 41789 && 
b[41790] == 41790 && 
b[41791] == 41791 && 
b[41792] == 41792 && 
b[41793] == 41793 && 
b[41794] == 41794 && 
b[41795] == 41795 && 
b[41796] == 41796 && 
b[41797] == 41797 && 
b[41798] == 41798 && 
b[41799] == 41799 && 
b[41800] == 41800 && 
b[41801] == 41801 && 
b[41802] == 41802 && 
b[41803] == 41803 && 
b[41804] == 41804 && 
b[41805] == 41805 && 
b[41806] == 41806 && 
b[41807] == 41807 && 
b[41808] == 41808 && 
b[41809] == 41809 && 
b[41810] == 41810 && 
b[41811] == 41811 && 
b[41812] == 41812 && 
b[41813] == 41813 && 
b[41814] == 41814 && 
b[41815] == 41815 && 
b[41816] == 41816 && 
b[41817] == 41817 && 
b[41818] == 41818 && 
b[41819] == 41819 && 
b[41820] == 41820 && 
b[41821] == 41821 && 
b[41822] == 41822 && 
b[41823] == 41823 && 
b[41824] == 41824 && 
b[41825] == 41825 && 
b[41826] == 41826 && 
b[41827] == 41827 && 
b[41828] == 41828 && 
b[41829] == 41829 && 
b[41830] == 41830 && 
b[41831] == 41831 && 
b[41832] == 41832 && 
b[41833] == 41833 && 
b[41834] == 41834 && 
b[41835] == 41835 && 
b[41836] == 41836 && 
b[41837] == 41837 && 
b[41838] == 41838 && 
b[41839] == 41839 && 
b[41840] == 41840 && 
b[41841] == 41841 && 
b[41842] == 41842 && 
b[41843] == 41843 && 
b[41844] == 41844 && 
b[41845] == 41845 && 
b[41846] == 41846 && 
b[41847] == 41847 && 
b[41848] == 41848 && 
b[41849] == 41849 && 
b[41850] == 41850 && 
b[41851] == 41851 && 
b[41852] == 41852 && 
b[41853] == 41853 && 
b[41854] == 41854 && 
b[41855] == 41855 && 
b[41856] == 41856 && 
b[41857] == 41857 && 
b[41858] == 41858 && 
b[41859] == 41859 && 
b[41860] == 41860 && 
b[41861] == 41861 && 
b[41862] == 41862 && 
b[41863] == 41863 && 
b[41864] == 41864 && 
b[41865] == 41865 && 
b[41866] == 41866 && 
b[41867] == 41867 && 
b[41868] == 41868 && 
b[41869] == 41869 && 
b[41870] == 41870 && 
b[41871] == 41871 && 
b[41872] == 41872 && 
b[41873] == 41873 && 
b[41874] == 41874 && 
b[41875] == 41875 && 
b[41876] == 41876 && 
b[41877] == 41877 && 
b[41878] == 41878 && 
b[41879] == 41879 && 
b[41880] == 41880 && 
b[41881] == 41881 && 
b[41882] == 41882 && 
b[41883] == 41883 && 
b[41884] == 41884 && 
b[41885] == 41885 && 
b[41886] == 41886 && 
b[41887] == 41887 && 
b[41888] == 41888 && 
b[41889] == 41889 && 
b[41890] == 41890 && 
b[41891] == 41891 && 
b[41892] == 41892 && 
b[41893] == 41893 && 
b[41894] == 41894 && 
b[41895] == 41895 && 
b[41896] == 41896 && 
b[41897] == 41897 && 
b[41898] == 41898 && 
b[41899] == 41899 && 
b[41900] == 41900 && 
b[41901] == 41901 && 
b[41902] == 41902 && 
b[41903] == 41903 && 
b[41904] == 41904 && 
b[41905] == 41905 && 
b[41906] == 41906 && 
b[41907] == 41907 && 
b[41908] == 41908 && 
b[41909] == 41909 && 
b[41910] == 41910 && 
b[41911] == 41911 && 
b[41912] == 41912 && 
b[41913] == 41913 && 
b[41914] == 41914 && 
b[41915] == 41915 && 
b[41916] == 41916 && 
b[41917] == 41917 && 
b[41918] == 41918 && 
b[41919] == 41919 && 
b[41920] == 41920 && 
b[41921] == 41921 && 
b[41922] == 41922 && 
b[41923] == 41923 && 
b[41924] == 41924 && 
b[41925] == 41925 && 
b[41926] == 41926 && 
b[41927] == 41927 && 
b[41928] == 41928 && 
b[41929] == 41929 && 
b[41930] == 41930 && 
b[41931] == 41931 && 
b[41932] == 41932 && 
b[41933] == 41933 && 
b[41934] == 41934 && 
b[41935] == 41935 && 
b[41936] == 41936 && 
b[41937] == 41937 && 
b[41938] == 41938 && 
b[41939] == 41939 && 
b[41940] == 41940 && 
b[41941] == 41941 && 
b[41942] == 41942 && 
b[41943] == 41943 && 
b[41944] == 41944 && 
b[41945] == 41945 && 
b[41946] == 41946 && 
b[41947] == 41947 && 
b[41948] == 41948 && 
b[41949] == 41949 && 
b[41950] == 41950 && 
b[41951] == 41951 && 
b[41952] == 41952 && 
b[41953] == 41953 && 
b[41954] == 41954 && 
b[41955] == 41955 && 
b[41956] == 41956 && 
b[41957] == 41957 && 
b[41958] == 41958 && 
b[41959] == 41959 && 
b[41960] == 41960 && 
b[41961] == 41961 && 
b[41962] == 41962 && 
b[41963] == 41963 && 
b[41964] == 41964 && 
b[41965] == 41965 && 
b[41966] == 41966 && 
b[41967] == 41967 && 
b[41968] == 41968 && 
b[41969] == 41969 && 
b[41970] == 41970 && 
b[41971] == 41971 && 
b[41972] == 41972 && 
b[41973] == 41973 && 
b[41974] == 41974 && 
b[41975] == 41975 && 
b[41976] == 41976 && 
b[41977] == 41977 && 
b[41978] == 41978 && 
b[41979] == 41979 && 
b[41980] == 41980 && 
b[41981] == 41981 && 
b[41982] == 41982 && 
b[41983] == 41983 && 
b[41984] == 41984 && 
b[41985] == 41985 && 
b[41986] == 41986 && 
b[41987] == 41987 && 
b[41988] == 41988 && 
b[41989] == 41989 && 
b[41990] == 41990 && 
b[41991] == 41991 && 
b[41992] == 41992 && 
b[41993] == 41993 && 
b[41994] == 41994 && 
b[41995] == 41995 && 
b[41996] == 41996 && 
b[41997] == 41997 && 
b[41998] == 41998 && 
b[41999] == 41999 && 
b[42000] == 42000 && 
b[42001] == 42001 && 
b[42002] == 42002 && 
b[42003] == 42003 && 
b[42004] == 42004 && 
b[42005] == 42005 && 
b[42006] == 42006 && 
b[42007] == 42007 && 
b[42008] == 42008 && 
b[42009] == 42009 && 
b[42010] == 42010 && 
b[42011] == 42011 && 
b[42012] == 42012 && 
b[42013] == 42013 && 
b[42014] == 42014 && 
b[42015] == 42015 && 
b[42016] == 42016 && 
b[42017] == 42017 && 
b[42018] == 42018 && 
b[42019] == 42019 && 
b[42020] == 42020 && 
b[42021] == 42021 && 
b[42022] == 42022 && 
b[42023] == 42023 && 
b[42024] == 42024 && 
b[42025] == 42025 && 
b[42026] == 42026 && 
b[42027] == 42027 && 
b[42028] == 42028 && 
b[42029] == 42029 && 
b[42030] == 42030 && 
b[42031] == 42031 && 
b[42032] == 42032 && 
b[42033] == 42033 && 
b[42034] == 42034 && 
b[42035] == 42035 && 
b[42036] == 42036 && 
b[42037] == 42037 && 
b[42038] == 42038 && 
b[42039] == 42039 && 
b[42040] == 42040 && 
b[42041] == 42041 && 
b[42042] == 42042 && 
b[42043] == 42043 && 
b[42044] == 42044 && 
b[42045] == 42045 && 
b[42046] == 42046 && 
b[42047] == 42047 && 
b[42048] == 42048 && 
b[42049] == 42049 && 
b[42050] == 42050 && 
b[42051] == 42051 && 
b[42052] == 42052 && 
b[42053] == 42053 && 
b[42054] == 42054 && 
b[42055] == 42055 && 
b[42056] == 42056 && 
b[42057] == 42057 && 
b[42058] == 42058 && 
b[42059] == 42059 && 
b[42060] == 42060 && 
b[42061] == 42061 && 
b[42062] == 42062 && 
b[42063] == 42063 && 
b[42064] == 42064 && 
b[42065] == 42065 && 
b[42066] == 42066 && 
b[42067] == 42067 && 
b[42068] == 42068 && 
b[42069] == 42069 && 
b[42070] == 42070 && 
b[42071] == 42071 && 
b[42072] == 42072 && 
b[42073] == 42073 && 
b[42074] == 42074 && 
b[42075] == 42075 && 
b[42076] == 42076 && 
b[42077] == 42077 && 
b[42078] == 42078 && 
b[42079] == 42079 && 
b[42080] == 42080 && 
b[42081] == 42081 && 
b[42082] == 42082 && 
b[42083] == 42083 && 
b[42084] == 42084 && 
b[42085] == 42085 && 
b[42086] == 42086 && 
b[42087] == 42087 && 
b[42088] == 42088 && 
b[42089] == 42089 && 
b[42090] == 42090 && 
b[42091] == 42091 && 
b[42092] == 42092 && 
b[42093] == 42093 && 
b[42094] == 42094 && 
b[42095] == 42095 && 
b[42096] == 42096 && 
b[42097] == 42097 && 
b[42098] == 42098 && 
b[42099] == 42099 && 
b[42100] == 42100 && 
b[42101] == 42101 && 
b[42102] == 42102 && 
b[42103] == 42103 && 
b[42104] == 42104 && 
b[42105] == 42105 && 
b[42106] == 42106 && 
b[42107] == 42107 && 
b[42108] == 42108 && 
b[42109] == 42109 && 
b[42110] == 42110 && 
b[42111] == 42111 && 
b[42112] == 42112 && 
b[42113] == 42113 && 
b[42114] == 42114 && 
b[42115] == 42115 && 
b[42116] == 42116 && 
b[42117] == 42117 && 
b[42118] == 42118 && 
b[42119] == 42119 && 
b[42120] == 42120 && 
b[42121] == 42121 && 
b[42122] == 42122 && 
b[42123] == 42123 && 
b[42124] == 42124 && 
b[42125] == 42125 && 
b[42126] == 42126 && 
b[42127] == 42127 && 
b[42128] == 42128 && 
b[42129] == 42129 && 
b[42130] == 42130 && 
b[42131] == 42131 && 
b[42132] == 42132 && 
b[42133] == 42133 && 
b[42134] == 42134 && 
b[42135] == 42135 && 
b[42136] == 42136 && 
b[42137] == 42137 && 
b[42138] == 42138 && 
b[42139] == 42139 && 
b[42140] == 42140 && 
b[42141] == 42141 && 
b[42142] == 42142 && 
b[42143] == 42143 && 
b[42144] == 42144 && 
b[42145] == 42145 && 
b[42146] == 42146 && 
b[42147] == 42147 && 
b[42148] == 42148 && 
b[42149] == 42149 && 
b[42150] == 42150 && 
b[42151] == 42151 && 
b[42152] == 42152 && 
b[42153] == 42153 && 
b[42154] == 42154 && 
b[42155] == 42155 && 
b[42156] == 42156 && 
b[42157] == 42157 && 
b[42158] == 42158 && 
b[42159] == 42159 && 
b[42160] == 42160 && 
b[42161] == 42161 && 
b[42162] == 42162 && 
b[42163] == 42163 && 
b[42164] == 42164 && 
b[42165] == 42165 && 
b[42166] == 42166 && 
b[42167] == 42167 && 
b[42168] == 42168 && 
b[42169] == 42169 && 
b[42170] == 42170 && 
b[42171] == 42171 && 
b[42172] == 42172 && 
b[42173] == 42173 && 
b[42174] == 42174 && 
b[42175] == 42175 && 
b[42176] == 42176 && 
b[42177] == 42177 && 
b[42178] == 42178 && 
b[42179] == 42179 && 
b[42180] == 42180 && 
b[42181] == 42181 && 
b[42182] == 42182 && 
b[42183] == 42183 && 
b[42184] == 42184 && 
b[42185] == 42185 && 
b[42186] == 42186 && 
b[42187] == 42187 && 
b[42188] == 42188 && 
b[42189] == 42189 && 
b[42190] == 42190 && 
b[42191] == 42191 && 
b[42192] == 42192 && 
b[42193] == 42193 && 
b[42194] == 42194 && 
b[42195] == 42195 && 
b[42196] == 42196 && 
b[42197] == 42197 && 
b[42198] == 42198 && 
b[42199] == 42199 && 
b[42200] == 42200 && 
b[42201] == 42201 && 
b[42202] == 42202 && 
b[42203] == 42203 && 
b[42204] == 42204 && 
b[42205] == 42205 && 
b[42206] == 42206 && 
b[42207] == 42207 && 
b[42208] == 42208 && 
b[42209] == 42209 && 
b[42210] == 42210 && 
b[42211] == 42211 && 
b[42212] == 42212 && 
b[42213] == 42213 && 
b[42214] == 42214 && 
b[42215] == 42215 && 
b[42216] == 42216 && 
b[42217] == 42217 && 
b[42218] == 42218 && 
b[42219] == 42219 && 
b[42220] == 42220 && 
b[42221] == 42221 && 
b[42222] == 42222 && 
b[42223] == 42223 && 
b[42224] == 42224 && 
b[42225] == 42225 && 
b[42226] == 42226 && 
b[42227] == 42227 && 
b[42228] == 42228 && 
b[42229] == 42229 && 
b[42230] == 42230 && 
b[42231] == 42231 && 
b[42232] == 42232 && 
b[42233] == 42233 && 
b[42234] == 42234 && 
b[42235] == 42235 && 
b[42236] == 42236 && 
b[42237] == 42237 && 
b[42238] == 42238 && 
b[42239] == 42239 && 
b[42240] == 42240 && 
b[42241] == 42241 && 
b[42242] == 42242 && 
b[42243] == 42243 && 
b[42244] == 42244 && 
b[42245] == 42245 && 
b[42246] == 42246 && 
b[42247] == 42247 && 
b[42248] == 42248 && 
b[42249] == 42249 && 
b[42250] == 42250 && 
b[42251] == 42251 && 
b[42252] == 42252 && 
b[42253] == 42253 && 
b[42254] == 42254 && 
b[42255] == 42255 && 
b[42256] == 42256 && 
b[42257] == 42257 && 
b[42258] == 42258 && 
b[42259] == 42259 && 
b[42260] == 42260 && 
b[42261] == 42261 && 
b[42262] == 42262 && 
b[42263] == 42263 && 
b[42264] == 42264 && 
b[42265] == 42265 && 
b[42266] == 42266 && 
b[42267] == 42267 && 
b[42268] == 42268 && 
b[42269] == 42269 && 
b[42270] == 42270 && 
b[42271] == 42271 && 
b[42272] == 42272 && 
b[42273] == 42273 && 
b[42274] == 42274 && 
b[42275] == 42275 && 
b[42276] == 42276 && 
b[42277] == 42277 && 
b[42278] == 42278 && 
b[42279] == 42279 && 
b[42280] == 42280 && 
b[42281] == 42281 && 
b[42282] == 42282 && 
b[42283] == 42283 && 
b[42284] == 42284 && 
b[42285] == 42285 && 
b[42286] == 42286 && 
b[42287] == 42287 && 
b[42288] == 42288 && 
b[42289] == 42289 && 
b[42290] == 42290 && 
b[42291] == 42291 && 
b[42292] == 42292 && 
b[42293] == 42293 && 
b[42294] == 42294 && 
b[42295] == 42295 && 
b[42296] == 42296 && 
b[42297] == 42297 && 
b[42298] == 42298 && 
b[42299] == 42299 && 
b[42300] == 42300 && 
b[42301] == 42301 && 
b[42302] == 42302 && 
b[42303] == 42303 && 
b[42304] == 42304 && 
b[42305] == 42305 && 
b[42306] == 42306 && 
b[42307] == 42307 && 
b[42308] == 42308 && 
b[42309] == 42309 && 
b[42310] == 42310 && 
b[42311] == 42311 && 
b[42312] == 42312 && 
b[42313] == 42313 && 
b[42314] == 42314 && 
b[42315] == 42315 && 
b[42316] == 42316 && 
b[42317] == 42317 && 
b[42318] == 42318 && 
b[42319] == 42319 && 
b[42320] == 42320 && 
b[42321] == 42321 && 
b[42322] == 42322 && 
b[42323] == 42323 && 
b[42324] == 42324 && 
b[42325] == 42325 && 
b[42326] == 42326 && 
b[42327] == 42327 && 
b[42328] == 42328 && 
b[42329] == 42329 && 
b[42330] == 42330 && 
b[42331] == 42331 && 
b[42332] == 42332 && 
b[42333] == 42333 && 
b[42334] == 42334 && 
b[42335] == 42335 && 
b[42336] == 42336 && 
b[42337] == 42337 && 
b[42338] == 42338 && 
b[42339] == 42339 && 
b[42340] == 42340 && 
b[42341] == 42341 && 
b[42342] == 42342 && 
b[42343] == 42343 && 
b[42344] == 42344 && 
b[42345] == 42345 && 
b[42346] == 42346 && 
b[42347] == 42347 && 
b[42348] == 42348 && 
b[42349] == 42349 && 
b[42350] == 42350 && 
b[42351] == 42351 && 
b[42352] == 42352 && 
b[42353] == 42353 && 
b[42354] == 42354 && 
b[42355] == 42355 && 
b[42356] == 42356 && 
b[42357] == 42357 && 
b[42358] == 42358 && 
b[42359] == 42359 && 
b[42360] == 42360 && 
b[42361] == 42361 && 
b[42362] == 42362 && 
b[42363] == 42363 && 
b[42364] == 42364 && 
b[42365] == 42365 && 
b[42366] == 42366 && 
b[42367] == 42367 && 
b[42368] == 42368 && 
b[42369] == 42369 && 
b[42370] == 42370 && 
b[42371] == 42371 && 
b[42372] == 42372 && 
b[42373] == 42373 && 
b[42374] == 42374 && 
b[42375] == 42375 && 
b[42376] == 42376 && 
b[42377] == 42377 && 
b[42378] == 42378 && 
b[42379] == 42379 && 
b[42380] == 42380 && 
b[42381] == 42381 && 
b[42382] == 42382 && 
b[42383] == 42383 && 
b[42384] == 42384 && 
b[42385] == 42385 && 
b[42386] == 42386 && 
b[42387] == 42387 && 
b[42388] == 42388 && 
b[42389] == 42389 && 
b[42390] == 42390 && 
b[42391] == 42391 && 
b[42392] == 42392 && 
b[42393] == 42393 && 
b[42394] == 42394 && 
b[42395] == 42395 && 
b[42396] == 42396 && 
b[42397] == 42397 && 
b[42398] == 42398 && 
b[42399] == 42399 && 
b[42400] == 42400 && 
b[42401] == 42401 && 
b[42402] == 42402 && 
b[42403] == 42403 && 
b[42404] == 42404 && 
b[42405] == 42405 && 
b[42406] == 42406 && 
b[42407] == 42407 && 
b[42408] == 42408 && 
b[42409] == 42409 && 
b[42410] == 42410 && 
b[42411] == 42411 && 
b[42412] == 42412 && 
b[42413] == 42413 && 
b[42414] == 42414 && 
b[42415] == 42415 && 
b[42416] == 42416 && 
b[42417] == 42417 && 
b[42418] == 42418 && 
b[42419] == 42419 && 
b[42420] == 42420 && 
b[42421] == 42421 && 
b[42422] == 42422 && 
b[42423] == 42423 && 
b[42424] == 42424 && 
b[42425] == 42425 && 
b[42426] == 42426 && 
b[42427] == 42427 && 
b[42428] == 42428 && 
b[42429] == 42429 && 
b[42430] == 42430 && 
b[42431] == 42431 && 
b[42432] == 42432 && 
b[42433] == 42433 && 
b[42434] == 42434 && 
b[42435] == 42435 && 
b[42436] == 42436 && 
b[42437] == 42437 && 
b[42438] == 42438 && 
b[42439] == 42439 && 
b[42440] == 42440 && 
b[42441] == 42441 && 
b[42442] == 42442 && 
b[42443] == 42443 && 
b[42444] == 42444 && 
b[42445] == 42445 && 
b[42446] == 42446 && 
b[42447] == 42447 && 
b[42448] == 42448 && 
b[42449] == 42449 && 
b[42450] == 42450 && 
b[42451] == 42451 && 
b[42452] == 42452 && 
b[42453] == 42453 && 
b[42454] == 42454 && 
b[42455] == 42455 && 
b[42456] == 42456 && 
b[42457] == 42457 && 
b[42458] == 42458 && 
b[42459] == 42459 && 
b[42460] == 42460 && 
b[42461] == 42461 && 
b[42462] == 42462 && 
b[42463] == 42463 && 
b[42464] == 42464 && 
b[42465] == 42465 && 
b[42466] == 42466 && 
b[42467] == 42467 && 
b[42468] == 42468 && 
b[42469] == 42469 && 
b[42470] == 42470 && 
b[42471] == 42471 && 
b[42472] == 42472 && 
b[42473] == 42473 && 
b[42474] == 42474 && 
b[42475] == 42475 && 
b[42476] == 42476 && 
b[42477] == 42477 && 
b[42478] == 42478 && 
b[42479] == 42479 && 
b[42480] == 42480 && 
b[42481] == 42481 && 
b[42482] == 42482 && 
b[42483] == 42483 && 
b[42484] == 42484 && 
b[42485] == 42485 && 
b[42486] == 42486 && 
b[42487] == 42487 && 
b[42488] == 42488 && 
b[42489] == 42489 && 
b[42490] == 42490 && 
b[42491] == 42491 && 
b[42492] == 42492 && 
b[42493] == 42493 && 
b[42494] == 42494 && 
b[42495] == 42495 && 
b[42496] == 42496 && 
b[42497] == 42497 && 
b[42498] == 42498 && 
b[42499] == 42499 && 
b[42500] == 42500 && 
b[42501] == 42501 && 
b[42502] == 42502 && 
b[42503] == 42503 && 
b[42504] == 42504 && 
b[42505] == 42505 && 
b[42506] == 42506 && 
b[42507] == 42507 && 
b[42508] == 42508 && 
b[42509] == 42509 && 
b[42510] == 42510 && 
b[42511] == 42511 && 
b[42512] == 42512 && 
b[42513] == 42513 && 
b[42514] == 42514 && 
b[42515] == 42515 && 
b[42516] == 42516 && 
b[42517] == 42517 && 
b[42518] == 42518 && 
b[42519] == 42519 && 
b[42520] == 42520 && 
b[42521] == 42521 && 
b[42522] == 42522 && 
b[42523] == 42523 && 
b[42524] == 42524 && 
b[42525] == 42525 && 
b[42526] == 42526 && 
b[42527] == 42527 && 
b[42528] == 42528 && 
b[42529] == 42529 && 
b[42530] == 42530 && 
b[42531] == 42531 && 
b[42532] == 42532 && 
b[42533] == 42533 && 
b[42534] == 42534 && 
b[42535] == 42535 && 
b[42536] == 42536 && 
b[42537] == 42537 && 
b[42538] == 42538 && 
b[42539] == 42539 && 
b[42540] == 42540 && 
b[42541] == 42541 && 
b[42542] == 42542 && 
b[42543] == 42543 && 
b[42544] == 42544 && 
b[42545] == 42545 && 
b[42546] == 42546 && 
b[42547] == 42547 && 
b[42548] == 42548 && 
b[42549] == 42549 && 
b[42550] == 42550 && 
b[42551] == 42551 && 
b[42552] == 42552 && 
b[42553] == 42553 && 
b[42554] == 42554 && 
b[42555] == 42555 && 
b[42556] == 42556 && 
b[42557] == 42557 && 
b[42558] == 42558 && 
b[42559] == 42559 && 
b[42560] == 42560 && 
b[42561] == 42561 && 
b[42562] == 42562 && 
b[42563] == 42563 && 
b[42564] == 42564 && 
b[42565] == 42565 && 
b[42566] == 42566 && 
b[42567] == 42567 && 
b[42568] == 42568 && 
b[42569] == 42569 && 
b[42570] == 42570 && 
b[42571] == 42571 && 
b[42572] == 42572 && 
b[42573] == 42573 && 
b[42574] == 42574 && 
b[42575] == 42575 && 
b[42576] == 42576 && 
b[42577] == 42577 && 
b[42578] == 42578 && 
b[42579] == 42579 && 
b[42580] == 42580 && 
b[42581] == 42581 && 
b[42582] == 42582 && 
b[42583] == 42583 && 
b[42584] == 42584 && 
b[42585] == 42585 && 
b[42586] == 42586 && 
b[42587] == 42587 && 
b[42588] == 42588 && 
b[42589] == 42589 && 
b[42590] == 42590 && 
b[42591] == 42591 && 
b[42592] == 42592 && 
b[42593] == 42593 && 
b[42594] == 42594 && 
b[42595] == 42595 && 
b[42596] == 42596 && 
b[42597] == 42597 && 
b[42598] == 42598 && 
b[42599] == 42599 && 
b[42600] == 42600 && 
b[42601] == 42601 && 
b[42602] == 42602 && 
b[42603] == 42603 && 
b[42604] == 42604 && 
b[42605] == 42605 && 
b[42606] == 42606 && 
b[42607] == 42607 && 
b[42608] == 42608 && 
b[42609] == 42609 && 
b[42610] == 42610 && 
b[42611] == 42611 && 
b[42612] == 42612 && 
b[42613] == 42613 && 
b[42614] == 42614 && 
b[42615] == 42615 && 
b[42616] == 42616 && 
b[42617] == 42617 && 
b[42618] == 42618 && 
b[42619] == 42619 && 
b[42620] == 42620 && 
b[42621] == 42621 && 
b[42622] == 42622 && 
b[42623] == 42623 && 
b[42624] == 42624 && 
b[42625] == 42625 && 
b[42626] == 42626 && 
b[42627] == 42627 && 
b[42628] == 42628 && 
b[42629] == 42629 && 
b[42630] == 42630 && 
b[42631] == 42631 && 
b[42632] == 42632 && 
b[42633] == 42633 && 
b[42634] == 42634 && 
b[42635] == 42635 && 
b[42636] == 42636 && 
b[42637] == 42637 && 
b[42638] == 42638 && 
b[42639] == 42639 && 
b[42640] == 42640 && 
b[42641] == 42641 && 
b[42642] == 42642 && 
b[42643] == 42643 && 
b[42644] == 42644 && 
b[42645] == 42645 && 
b[42646] == 42646 && 
b[42647] == 42647 && 
b[42648] == 42648 && 
b[42649] == 42649 && 
b[42650] == 42650 && 
b[42651] == 42651 && 
b[42652] == 42652 && 
b[42653] == 42653 && 
b[42654] == 42654 && 
b[42655] == 42655 && 
b[42656] == 42656 && 
b[42657] == 42657 && 
b[42658] == 42658 && 
b[42659] == 42659 && 
b[42660] == 42660 && 
b[42661] == 42661 && 
b[42662] == 42662 && 
b[42663] == 42663 && 
b[42664] == 42664 && 
b[42665] == 42665 && 
b[42666] == 42666 && 
b[42667] == 42667 && 
b[42668] == 42668 && 
b[42669] == 42669 && 
b[42670] == 42670 && 
b[42671] == 42671 && 
b[42672] == 42672 && 
b[42673] == 42673 && 
b[42674] == 42674 && 
b[42675] == 42675 && 
b[42676] == 42676 && 
b[42677] == 42677 && 
b[42678] == 42678 && 
b[42679] == 42679 && 
b[42680] == 42680 && 
b[42681] == 42681 && 
b[42682] == 42682 && 
b[42683] == 42683 && 
b[42684] == 42684 && 
b[42685] == 42685 && 
b[42686] == 42686 && 
b[42687] == 42687 && 
b[42688] == 42688 && 
b[42689] == 42689 && 
b[42690] == 42690 && 
b[42691] == 42691 && 
b[42692] == 42692 && 
b[42693] == 42693 && 
b[42694] == 42694 && 
b[42695] == 42695 && 
b[42696] == 42696 && 
b[42697] == 42697 && 
b[42698] == 42698 && 
b[42699] == 42699 && 
b[42700] == 42700 && 
b[42701] == 42701 && 
b[42702] == 42702 && 
b[42703] == 42703 && 
b[42704] == 42704 && 
b[42705] == 42705 && 
b[42706] == 42706 && 
b[42707] == 42707 && 
b[42708] == 42708 && 
b[42709] == 42709 && 
b[42710] == 42710 && 
b[42711] == 42711 && 
b[42712] == 42712 && 
b[42713] == 42713 && 
b[42714] == 42714 && 
b[42715] == 42715 && 
b[42716] == 42716 && 
b[42717] == 42717 && 
b[42718] == 42718 && 
b[42719] == 42719 && 
b[42720] == 42720 && 
b[42721] == 42721 && 
b[42722] == 42722 && 
b[42723] == 42723 && 
b[42724] == 42724 && 
b[42725] == 42725 && 
b[42726] == 42726 && 
b[42727] == 42727 && 
b[42728] == 42728 && 
b[42729] == 42729 && 
b[42730] == 42730 && 
b[42731] == 42731 && 
b[42732] == 42732 && 
b[42733] == 42733 && 
b[42734] == 42734 && 
b[42735] == 42735 && 
b[42736] == 42736 && 
b[42737] == 42737 && 
b[42738] == 42738 && 
b[42739] == 42739 && 
b[42740] == 42740 && 
b[42741] == 42741 && 
b[42742] == 42742 && 
b[42743] == 42743 && 
b[42744] == 42744 && 
b[42745] == 42745 && 
b[42746] == 42746 && 
b[42747] == 42747 && 
b[42748] == 42748 && 
b[42749] == 42749 && 
b[42750] == 42750 && 
b[42751] == 42751 && 
b[42752] == 42752 && 
b[42753] == 42753 && 
b[42754] == 42754 && 
b[42755] == 42755 && 
b[42756] == 42756 && 
b[42757] == 42757 && 
b[42758] == 42758 && 
b[42759] == 42759 && 
b[42760] == 42760 && 
b[42761] == 42761 && 
b[42762] == 42762 && 
b[42763] == 42763 && 
b[42764] == 42764 && 
b[42765] == 42765 && 
b[42766] == 42766 && 
b[42767] == 42767 && 
b[42768] == 42768 && 
b[42769] == 42769 && 
b[42770] == 42770 && 
b[42771] == 42771 && 
b[42772] == 42772 && 
b[42773] == 42773 && 
b[42774] == 42774 && 
b[42775] == 42775 && 
b[42776] == 42776 && 
b[42777] == 42777 && 
b[42778] == 42778 && 
b[42779] == 42779 && 
b[42780] == 42780 && 
b[42781] == 42781 && 
b[42782] == 42782 && 
b[42783] == 42783 && 
b[42784] == 42784 && 
b[42785] == 42785 && 
b[42786] == 42786 && 
b[42787] == 42787 && 
b[42788] == 42788 && 
b[42789] == 42789 && 
b[42790] == 42790 && 
b[42791] == 42791 && 
b[42792] == 42792 && 
b[42793] == 42793 && 
b[42794] == 42794 && 
b[42795] == 42795 && 
b[42796] == 42796 && 
b[42797] == 42797 && 
b[42798] == 42798 && 
b[42799] == 42799 && 
b[42800] == 42800 && 
b[42801] == 42801 && 
b[42802] == 42802 && 
b[42803] == 42803 && 
b[42804] == 42804 && 
b[42805] == 42805 && 
b[42806] == 42806 && 
b[42807] == 42807 && 
b[42808] == 42808 && 
b[42809] == 42809 && 
b[42810] == 42810 && 
b[42811] == 42811 && 
b[42812] == 42812 && 
b[42813] == 42813 && 
b[42814] == 42814 && 
b[42815] == 42815 && 
b[42816] == 42816 && 
b[42817] == 42817 && 
b[42818] == 42818 && 
b[42819] == 42819 && 
b[42820] == 42820 && 
b[42821] == 42821 && 
b[42822] == 42822 && 
b[42823] == 42823 && 
b[42824] == 42824 && 
b[42825] == 42825 && 
b[42826] == 42826 && 
b[42827] == 42827 && 
b[42828] == 42828 && 
b[42829] == 42829 && 
b[42830] == 42830 && 
b[42831] == 42831 && 
b[42832] == 42832 && 
b[42833] == 42833 && 
b[42834] == 42834 && 
b[42835] == 42835 && 
b[42836] == 42836 && 
b[42837] == 42837 && 
b[42838] == 42838 && 
b[42839] == 42839 && 
b[42840] == 42840 && 
b[42841] == 42841 && 
b[42842] == 42842 && 
b[42843] == 42843 && 
b[42844] == 42844 && 
b[42845] == 42845 && 
b[42846] == 42846 && 
b[42847] == 42847 && 
b[42848] == 42848 && 
b[42849] == 42849 && 
b[42850] == 42850 && 
b[42851] == 42851 && 
b[42852] == 42852 && 
b[42853] == 42853 && 
b[42854] == 42854 && 
b[42855] == 42855 && 
b[42856] == 42856 && 
b[42857] == 42857 && 
b[42858] == 42858 && 
b[42859] == 42859 && 
b[42860] == 42860 && 
b[42861] == 42861 && 
b[42862] == 42862 && 
b[42863] == 42863 && 
b[42864] == 42864 && 
b[42865] == 42865 && 
b[42866] == 42866 && 
b[42867] == 42867 && 
b[42868] == 42868 && 
b[42869] == 42869 && 
b[42870] == 42870 && 
b[42871] == 42871 && 
b[42872] == 42872 && 
b[42873] == 42873 && 
b[42874] == 42874 && 
b[42875] == 42875 && 
b[42876] == 42876 && 
b[42877] == 42877 && 
b[42878] == 42878 && 
b[42879] == 42879 && 
b[42880] == 42880 && 
b[42881] == 42881 && 
b[42882] == 42882 && 
b[42883] == 42883 && 
b[42884] == 42884 && 
b[42885] == 42885 && 
b[42886] == 42886 && 
b[42887] == 42887 && 
b[42888] == 42888 && 
b[42889] == 42889 && 
b[42890] == 42890 && 
b[42891] == 42891 && 
b[42892] == 42892 && 
b[42893] == 42893 && 
b[42894] == 42894 && 
b[42895] == 42895 && 
b[42896] == 42896 && 
b[42897] == 42897 && 
b[42898] == 42898 && 
b[42899] == 42899 && 
b[42900] == 42900 && 
b[42901] == 42901 && 
b[42902] == 42902 && 
b[42903] == 42903 && 
b[42904] == 42904 && 
b[42905] == 42905 && 
b[42906] == 42906 && 
b[42907] == 42907 && 
b[42908] == 42908 && 
b[42909] == 42909 && 
b[42910] == 42910 && 
b[42911] == 42911 && 
b[42912] == 42912 && 
b[42913] == 42913 && 
b[42914] == 42914 && 
b[42915] == 42915 && 
b[42916] == 42916 && 
b[42917] == 42917 && 
b[42918] == 42918 && 
b[42919] == 42919 && 
b[42920] == 42920 && 
b[42921] == 42921 && 
b[42922] == 42922 && 
b[42923] == 42923 && 
b[42924] == 42924 && 
b[42925] == 42925 && 
b[42926] == 42926 && 
b[42927] == 42927 && 
b[42928] == 42928 && 
b[42929] == 42929 && 
b[42930] == 42930 && 
b[42931] == 42931 && 
b[42932] == 42932 && 
b[42933] == 42933 && 
b[42934] == 42934 && 
b[42935] == 42935 && 
b[42936] == 42936 && 
b[42937] == 42937 && 
b[42938] == 42938 && 
b[42939] == 42939 && 
b[42940] == 42940 && 
b[42941] == 42941 && 
b[42942] == 42942 && 
b[42943] == 42943 && 
b[42944] == 42944 && 
b[42945] == 42945 && 
b[42946] == 42946 && 
b[42947] == 42947 && 
b[42948] == 42948 && 
b[42949] == 42949 && 
b[42950] == 42950 && 
b[42951] == 42951 && 
b[42952] == 42952 && 
b[42953] == 42953 && 
b[42954] == 42954 && 
b[42955] == 42955 && 
b[42956] == 42956 && 
b[42957] == 42957 && 
b[42958] == 42958 && 
b[42959] == 42959 && 
b[42960] == 42960 && 
b[42961] == 42961 && 
b[42962] == 42962 && 
b[42963] == 42963 && 
b[42964] == 42964 && 
b[42965] == 42965 && 
b[42966] == 42966 && 
b[42967] == 42967 && 
b[42968] == 42968 && 
b[42969] == 42969 && 
b[42970] == 42970 && 
b[42971] == 42971 && 
b[42972] == 42972 && 
b[42973] == 42973 && 
b[42974] == 42974 && 
b[42975] == 42975 && 
b[42976] == 42976 && 
b[42977] == 42977 && 
b[42978] == 42978 && 
b[42979] == 42979 && 
b[42980] == 42980 && 
b[42981] == 42981 && 
b[42982] == 42982 && 
b[42983] == 42983 && 
b[42984] == 42984 && 
b[42985] == 42985 && 
b[42986] == 42986 && 
b[42987] == 42987 && 
b[42988] == 42988 && 
b[42989] == 42989 && 
b[42990] == 42990 && 
b[42991] == 42991 && 
b[42992] == 42992 && 
b[42993] == 42993 && 
b[42994] == 42994 && 
b[42995] == 42995 && 
b[42996] == 42996 && 
b[42997] == 42997 && 
b[42998] == 42998 && 
b[42999] == 42999 && 
b[43000] == 43000 && 
b[43001] == 43001 && 
b[43002] == 43002 && 
b[43003] == 43003 && 
b[43004] == 43004 && 
b[43005] == 43005 && 
b[43006] == 43006 && 
b[43007] == 43007 && 
b[43008] == 43008 && 
b[43009] == 43009 && 
b[43010] == 43010 && 
b[43011] == 43011 && 
b[43012] == 43012 && 
b[43013] == 43013 && 
b[43014] == 43014 && 
b[43015] == 43015 && 
b[43016] == 43016 && 
b[43017] == 43017 && 
b[43018] == 43018 && 
b[43019] == 43019 && 
b[43020] == 43020 && 
b[43021] == 43021 && 
b[43022] == 43022 && 
b[43023] == 43023 && 
b[43024] == 43024 && 
b[43025] == 43025 && 
b[43026] == 43026 && 
b[43027] == 43027 && 
b[43028] == 43028 && 
b[43029] == 43029 && 
b[43030] == 43030 && 
b[43031] == 43031 && 
b[43032] == 43032 && 
b[43033] == 43033 && 
b[43034] == 43034 && 
b[43035] == 43035 && 
b[43036] == 43036 && 
b[43037] == 43037 && 
b[43038] == 43038 && 
b[43039] == 43039 && 
b[43040] == 43040 && 
b[43041] == 43041 && 
b[43042] == 43042 && 
b[43043] == 43043 && 
b[43044] == 43044 && 
b[43045] == 43045 && 
b[43046] == 43046 && 
b[43047] == 43047 && 
b[43048] == 43048 && 
b[43049] == 43049 && 
b[43050] == 43050 && 
b[43051] == 43051 && 
b[43052] == 43052 && 
b[43053] == 43053 && 
b[43054] == 43054 && 
b[43055] == 43055 && 
b[43056] == 43056 && 
b[43057] == 43057 && 
b[43058] == 43058 && 
b[43059] == 43059 && 
b[43060] == 43060 && 
b[43061] == 43061 && 
b[43062] == 43062 && 
b[43063] == 43063 && 
b[43064] == 43064 && 
b[43065] == 43065 && 
b[43066] == 43066 && 
b[43067] == 43067 && 
b[43068] == 43068 && 
b[43069] == 43069 && 
b[43070] == 43070 && 
b[43071] == 43071 && 
b[43072] == 43072 && 
b[43073] == 43073 && 
b[43074] == 43074 && 
b[43075] == 43075 && 
b[43076] == 43076 && 
b[43077] == 43077 && 
b[43078] == 43078 && 
b[43079] == 43079 && 
b[43080] == 43080 && 
b[43081] == 43081 && 
b[43082] == 43082 && 
b[43083] == 43083 && 
b[43084] == 43084 && 
b[43085] == 43085 && 
b[43086] == 43086 && 
b[43087] == 43087 && 
b[43088] == 43088 && 
b[43089] == 43089 && 
b[43090] == 43090 && 
b[43091] == 43091 && 
b[43092] == 43092 && 
b[43093] == 43093 && 
b[43094] == 43094 && 
b[43095] == 43095 && 
b[43096] == 43096 && 
b[43097] == 43097 && 
b[43098] == 43098 && 
b[43099] == 43099 && 
b[43100] == 43100 && 
b[43101] == 43101 && 
b[43102] == 43102 && 
b[43103] == 43103 && 
b[43104] == 43104 && 
b[43105] == 43105 && 
b[43106] == 43106 && 
b[43107] == 43107 && 
b[43108] == 43108 && 
b[43109] == 43109 && 
b[43110] == 43110 && 
b[43111] == 43111 && 
b[43112] == 43112 && 
b[43113] == 43113 && 
b[43114] == 43114 && 
b[43115] == 43115 && 
b[43116] == 43116 && 
b[43117] == 43117 && 
b[43118] == 43118 && 
b[43119] == 43119 && 
b[43120] == 43120 && 
b[43121] == 43121 && 
b[43122] == 43122 && 
b[43123] == 43123 && 
b[43124] == 43124 && 
b[43125] == 43125 && 
b[43126] == 43126 && 
b[43127] == 43127 && 
b[43128] == 43128 && 
b[43129] == 43129 && 
b[43130] == 43130 && 
b[43131] == 43131 && 
b[43132] == 43132 && 
b[43133] == 43133 && 
b[43134] == 43134 && 
b[43135] == 43135 && 
b[43136] == 43136 && 
b[43137] == 43137 && 
b[43138] == 43138 && 
b[43139] == 43139 && 
b[43140] == 43140 && 
b[43141] == 43141 && 
b[43142] == 43142 && 
b[43143] == 43143 && 
b[43144] == 43144 && 
b[43145] == 43145 && 
b[43146] == 43146 && 
b[43147] == 43147 && 
b[43148] == 43148 && 
b[43149] == 43149 && 
b[43150] == 43150 && 
b[43151] == 43151 && 
b[43152] == 43152 && 
b[43153] == 43153 && 
b[43154] == 43154 && 
b[43155] == 43155 && 
b[43156] == 43156 && 
b[43157] == 43157 && 
b[43158] == 43158 && 
b[43159] == 43159 && 
b[43160] == 43160 && 
b[43161] == 43161 && 
b[43162] == 43162 && 
b[43163] == 43163 && 
b[43164] == 43164 && 
b[43165] == 43165 && 
b[43166] == 43166 && 
b[43167] == 43167 && 
b[43168] == 43168 && 
b[43169] == 43169 && 
b[43170] == 43170 && 
b[43171] == 43171 && 
b[43172] == 43172 && 
b[43173] == 43173 && 
b[43174] == 43174 && 
b[43175] == 43175 && 
b[43176] == 43176 && 
b[43177] == 43177 && 
b[43178] == 43178 && 
b[43179] == 43179 && 
b[43180] == 43180 && 
b[43181] == 43181 && 
b[43182] == 43182 && 
b[43183] == 43183 && 
b[43184] == 43184 && 
b[43185] == 43185 && 
b[43186] == 43186 && 
b[43187] == 43187 && 
b[43188] == 43188 && 
b[43189] == 43189 && 
b[43190] == 43190 && 
b[43191] == 43191 && 
b[43192] == 43192 && 
b[43193] == 43193 && 
b[43194] == 43194 && 
b[43195] == 43195 && 
b[43196] == 43196 && 
b[43197] == 43197 && 
b[43198] == 43198 && 
b[43199] == 43199 && 
b[43200] == 43200 && 
b[43201] == 43201 && 
b[43202] == 43202 && 
b[43203] == 43203 && 
b[43204] == 43204 && 
b[43205] == 43205 && 
b[43206] == 43206 && 
b[43207] == 43207 && 
b[43208] == 43208 && 
b[43209] == 43209 && 
b[43210] == 43210 && 
b[43211] == 43211 && 
b[43212] == 43212 && 
b[43213] == 43213 && 
b[43214] == 43214 && 
b[43215] == 43215 && 
b[43216] == 43216 && 
b[43217] == 43217 && 
b[43218] == 43218 && 
b[43219] == 43219 && 
b[43220] == 43220 && 
b[43221] == 43221 && 
b[43222] == 43222 && 
b[43223] == 43223 && 
b[43224] == 43224 && 
b[43225] == 43225 && 
b[43226] == 43226 && 
b[43227] == 43227 && 
b[43228] == 43228 && 
b[43229] == 43229 && 
b[43230] == 43230 && 
b[43231] == 43231 && 
b[43232] == 43232 && 
b[43233] == 43233 && 
b[43234] == 43234 && 
b[43235] == 43235 && 
b[43236] == 43236 && 
b[43237] == 43237 && 
b[43238] == 43238 && 
b[43239] == 43239 && 
b[43240] == 43240 && 
b[43241] == 43241 && 
b[43242] == 43242 && 
b[43243] == 43243 && 
b[43244] == 43244 && 
b[43245] == 43245 && 
b[43246] == 43246 && 
b[43247] == 43247 && 
b[43248] == 43248 && 
b[43249] == 43249 && 
b[43250] == 43250 && 
b[43251] == 43251 && 
b[43252] == 43252 && 
b[43253] == 43253 && 
b[43254] == 43254 && 
b[43255] == 43255 && 
b[43256] == 43256 && 
b[43257] == 43257 && 
b[43258] == 43258 && 
b[43259] == 43259 && 
b[43260] == 43260 && 
b[43261] == 43261 && 
b[43262] == 43262 && 
b[43263] == 43263 && 
b[43264] == 43264 && 
b[43265] == 43265 && 
b[43266] == 43266 && 
b[43267] == 43267 && 
b[43268] == 43268 && 
b[43269] == 43269 && 
b[43270] == 43270 && 
b[43271] == 43271 && 
b[43272] == 43272 && 
b[43273] == 43273 && 
b[43274] == 43274 && 
b[43275] == 43275 && 
b[43276] == 43276 && 
b[43277] == 43277 && 
b[43278] == 43278 && 
b[43279] == 43279 && 
b[43280] == 43280 && 
b[43281] == 43281 && 
b[43282] == 43282 && 
b[43283] == 43283 && 
b[43284] == 43284 && 
b[43285] == 43285 && 
b[43286] == 43286 && 
b[43287] == 43287 && 
b[43288] == 43288 && 
b[43289] == 43289 && 
b[43290] == 43290 && 
b[43291] == 43291 && 
b[43292] == 43292 && 
b[43293] == 43293 && 
b[43294] == 43294 && 
b[43295] == 43295 && 
b[43296] == 43296 && 
b[43297] == 43297 && 
b[43298] == 43298 && 
b[43299] == 43299 && 
b[43300] == 43300 && 
b[43301] == 43301 && 
b[43302] == 43302 && 
b[43303] == 43303 && 
b[43304] == 43304 && 
b[43305] == 43305 && 
b[43306] == 43306 && 
b[43307] == 43307 && 
b[43308] == 43308 && 
b[43309] == 43309 && 
b[43310] == 43310 && 
b[43311] == 43311 && 
b[43312] == 43312 && 
b[43313] == 43313 && 
b[43314] == 43314 && 
b[43315] == 43315 && 
b[43316] == 43316 && 
b[43317] == 43317 && 
b[43318] == 43318 && 
b[43319] == 43319 && 
b[43320] == 43320 && 
b[43321] == 43321 && 
b[43322] == 43322 && 
b[43323] == 43323 && 
b[43324] == 43324 && 
b[43325] == 43325 && 
b[43326] == 43326 && 
b[43327] == 43327 && 
b[43328] == 43328 && 
b[43329] == 43329 && 
b[43330] == 43330 && 
b[43331] == 43331 && 
b[43332] == 43332 && 
b[43333] == 43333 && 
b[43334] == 43334 && 
b[43335] == 43335 && 
b[43336] == 43336 && 
b[43337] == 43337 && 
b[43338] == 43338 && 
b[43339] == 43339 && 
b[43340] == 43340 && 
b[43341] == 43341 && 
b[43342] == 43342 && 
b[43343] == 43343 && 
b[43344] == 43344 && 
b[43345] == 43345 && 
b[43346] == 43346 && 
b[43347] == 43347 && 
b[43348] == 43348 && 
b[43349] == 43349 && 
b[43350] == 43350 && 
b[43351] == 43351 && 
b[43352] == 43352 && 
b[43353] == 43353 && 
b[43354] == 43354 && 
b[43355] == 43355 && 
b[43356] == 43356 && 
b[43357] == 43357 && 
b[43358] == 43358 && 
b[43359] == 43359 && 
b[43360] == 43360 && 
b[43361] == 43361 && 
b[43362] == 43362 && 
b[43363] == 43363 && 
b[43364] == 43364 && 
b[43365] == 43365 && 
b[43366] == 43366 && 
b[43367] == 43367 && 
b[43368] == 43368 && 
b[43369] == 43369 && 
b[43370] == 43370 && 
b[43371] == 43371 && 
b[43372] == 43372 && 
b[43373] == 43373 && 
b[43374] == 43374 && 
b[43375] == 43375 && 
b[43376] == 43376 && 
b[43377] == 43377 && 
b[43378] == 43378 && 
b[43379] == 43379 && 
b[43380] == 43380 && 
b[43381] == 43381 && 
b[43382] == 43382 && 
b[43383] == 43383 && 
b[43384] == 43384 && 
b[43385] == 43385 && 
b[43386] == 43386 && 
b[43387] == 43387 && 
b[43388] == 43388 && 
b[43389] == 43389 && 
b[43390] == 43390 && 
b[43391] == 43391 && 
b[43392] == 43392 && 
b[43393] == 43393 && 
b[43394] == 43394 && 
b[43395] == 43395 && 
b[43396] == 43396 && 
b[43397] == 43397 && 
b[43398] == 43398 && 
b[43399] == 43399 && 
b[43400] == 43400 && 
b[43401] == 43401 && 
b[43402] == 43402 && 
b[43403] == 43403 && 
b[43404] == 43404 && 
b[43405] == 43405 && 
b[43406] == 43406 && 
b[43407] == 43407 && 
b[43408] == 43408 && 
b[43409] == 43409 && 
b[43410] == 43410 && 
b[43411] == 43411 && 
b[43412] == 43412 && 
b[43413] == 43413 && 
b[43414] == 43414 && 
b[43415] == 43415 && 
b[43416] == 43416 && 
b[43417] == 43417 && 
b[43418] == 43418 && 
b[43419] == 43419 && 
b[43420] == 43420 && 
b[43421] == 43421 && 
b[43422] == 43422 && 
b[43423] == 43423 && 
b[43424] == 43424 && 
b[43425] == 43425 && 
b[43426] == 43426 && 
b[43427] == 43427 && 
b[43428] == 43428 && 
b[43429] == 43429 && 
b[43430] == 43430 && 
b[43431] == 43431 && 
b[43432] == 43432 && 
b[43433] == 43433 && 
b[43434] == 43434 && 
b[43435] == 43435 && 
b[43436] == 43436 && 
b[43437] == 43437 && 
b[43438] == 43438 && 
b[43439] == 43439 && 
b[43440] == 43440 && 
b[43441] == 43441 && 
b[43442] == 43442 && 
b[43443] == 43443 && 
b[43444] == 43444 && 
b[43445] == 43445 && 
b[43446] == 43446 && 
b[43447] == 43447 && 
b[43448] == 43448 && 
b[43449] == 43449 && 
b[43450] == 43450 && 
b[43451] == 43451 && 
b[43452] == 43452 && 
b[43453] == 43453 && 
b[43454] == 43454 && 
b[43455] == 43455 && 
b[43456] == 43456 && 
b[43457] == 43457 && 
b[43458] == 43458 && 
b[43459] == 43459 && 
b[43460] == 43460 && 
b[43461] == 43461 && 
b[43462] == 43462 && 
b[43463] == 43463 && 
b[43464] == 43464 && 
b[43465] == 43465 && 
b[43466] == 43466 && 
b[43467] == 43467 && 
b[43468] == 43468 && 
b[43469] == 43469 && 
b[43470] == 43470 && 
b[43471] == 43471 && 
b[43472] == 43472 && 
b[43473] == 43473 && 
b[43474] == 43474 && 
b[43475] == 43475 && 
b[43476] == 43476 && 
b[43477] == 43477 && 
b[43478] == 43478 && 
b[43479] == 43479 && 
b[43480] == 43480 && 
b[43481] == 43481 && 
b[43482] == 43482 && 
b[43483] == 43483 && 
b[43484] == 43484 && 
b[43485] == 43485 && 
b[43486] == 43486 && 
b[43487] == 43487 && 
b[43488] == 43488 && 
b[43489] == 43489 && 
b[43490] == 43490 && 
b[43491] == 43491 && 
b[43492] == 43492 && 
b[43493] == 43493 && 
b[43494] == 43494 && 
b[43495] == 43495 && 
b[43496] == 43496 && 
b[43497] == 43497 && 
b[43498] == 43498 && 
b[43499] == 43499 && 
b[43500] == 43500 && 
b[43501] == 43501 && 
b[43502] == 43502 && 
b[43503] == 43503 && 
b[43504] == 43504 && 
b[43505] == 43505 && 
b[43506] == 43506 && 
b[43507] == 43507 && 
b[43508] == 43508 && 
b[43509] == 43509 && 
b[43510] == 43510 && 
b[43511] == 43511 && 
b[43512] == 43512 && 
b[43513] == 43513 && 
b[43514] == 43514 && 
b[43515] == 43515 && 
b[43516] == 43516 && 
b[43517] == 43517 && 
b[43518] == 43518 && 
b[43519] == 43519 && 
b[43520] == 43520 && 
b[43521] == 43521 && 
b[43522] == 43522 && 
b[43523] == 43523 && 
b[43524] == 43524 && 
b[43525] == 43525 && 
b[43526] == 43526 && 
b[43527] == 43527 && 
b[43528] == 43528 && 
b[43529] == 43529 && 
b[43530] == 43530 && 
b[43531] == 43531 && 
b[43532] == 43532 && 
b[43533] == 43533 && 
b[43534] == 43534 && 
b[43535] == 43535 && 
b[43536] == 43536 && 
b[43537] == 43537 && 
b[43538] == 43538 && 
b[43539] == 43539 && 
b[43540] == 43540 && 
b[43541] == 43541 && 
b[43542] == 43542 && 
b[43543] == 43543 && 
b[43544] == 43544 && 
b[43545] == 43545 && 
b[43546] == 43546 && 
b[43547] == 43547 && 
b[43548] == 43548 && 
b[43549] == 43549 && 
b[43550] == 43550 && 
b[43551] == 43551 && 
b[43552] == 43552 && 
b[43553] == 43553 && 
b[43554] == 43554 && 
b[43555] == 43555 && 
b[43556] == 43556 && 
b[43557] == 43557 && 
b[43558] == 43558 && 
b[43559] == 43559 && 
b[43560] == 43560 && 
b[43561] == 43561 && 
b[43562] == 43562 && 
b[43563] == 43563 && 
b[43564] == 43564 && 
b[43565] == 43565 && 
b[43566] == 43566 && 
b[43567] == 43567 && 
b[43568] == 43568 && 
b[43569] == 43569 && 
b[43570] == 43570 && 
b[43571] == 43571 && 
b[43572] == 43572 && 
b[43573] == 43573 && 
b[43574] == 43574 && 
b[43575] == 43575 && 
b[43576] == 43576 && 
b[43577] == 43577 && 
b[43578] == 43578 && 
b[43579] == 43579 && 
b[43580] == 43580 && 
b[43581] == 43581 && 
b[43582] == 43582 && 
b[43583] == 43583 && 
b[43584] == 43584 && 
b[43585] == 43585 && 
b[43586] == 43586 && 
b[43587] == 43587 && 
b[43588] == 43588 && 
b[43589] == 43589 && 
b[43590] == 43590 && 
b[43591] == 43591 && 
b[43592] == 43592 && 
b[43593] == 43593 && 
b[43594] == 43594 && 
b[43595] == 43595 && 
b[43596] == 43596 && 
b[43597] == 43597 && 
b[43598] == 43598 && 
b[43599] == 43599 && 
b[43600] == 43600 && 
b[43601] == 43601 && 
b[43602] == 43602 && 
b[43603] == 43603 && 
b[43604] == 43604 && 
b[43605] == 43605 && 
b[43606] == 43606 && 
b[43607] == 43607 && 
b[43608] == 43608 && 
b[43609] == 43609 && 
b[43610] == 43610 && 
b[43611] == 43611 && 
b[43612] == 43612 && 
b[43613] == 43613 && 
b[43614] == 43614 && 
b[43615] == 43615 && 
b[43616] == 43616 && 
b[43617] == 43617 && 
b[43618] == 43618 && 
b[43619] == 43619 && 
b[43620] == 43620 && 
b[43621] == 43621 && 
b[43622] == 43622 && 
b[43623] == 43623 && 
b[43624] == 43624 && 
b[43625] == 43625 && 
b[43626] == 43626 && 
b[43627] == 43627 && 
b[43628] == 43628 && 
b[43629] == 43629 && 
b[43630] == 43630 && 
b[43631] == 43631 && 
b[43632] == 43632 && 
b[43633] == 43633 && 
b[43634] == 43634 && 
b[43635] == 43635 && 
b[43636] == 43636 && 
b[43637] == 43637 && 
b[43638] == 43638 && 
b[43639] == 43639 && 
b[43640] == 43640 && 
b[43641] == 43641 && 
b[43642] == 43642 && 
b[43643] == 43643 && 
b[43644] == 43644 && 
b[43645] == 43645 && 
b[43646] == 43646 && 
b[43647] == 43647 && 
b[43648] == 43648 && 
b[43649] == 43649 && 
b[43650] == 43650 && 
b[43651] == 43651 && 
b[43652] == 43652 && 
b[43653] == 43653 && 
b[43654] == 43654 && 
b[43655] == 43655 && 
b[43656] == 43656 && 
b[43657] == 43657 && 
b[43658] == 43658 && 
b[43659] == 43659 && 
b[43660] == 43660 && 
b[43661] == 43661 && 
b[43662] == 43662 && 
b[43663] == 43663 && 
b[43664] == 43664 && 
b[43665] == 43665 && 
b[43666] == 43666 && 
b[43667] == 43667 && 
b[43668] == 43668 && 
b[43669] == 43669 && 
b[43670] == 43670 && 
b[43671] == 43671 && 
b[43672] == 43672 && 
b[43673] == 43673 && 
b[43674] == 43674 && 
b[43675] == 43675 && 
b[43676] == 43676 && 
b[43677] == 43677 && 
b[43678] == 43678 && 
b[43679] == 43679 && 
b[43680] == 43680 && 
b[43681] == 43681 && 
b[43682] == 43682 && 
b[43683] == 43683 && 
b[43684] == 43684 && 
b[43685] == 43685 && 
b[43686] == 43686 && 
b[43687] == 43687 && 
b[43688] == 43688 && 
b[43689] == 43689 && 
b[43690] == 43690 && 
b[43691] == 43691 && 
b[43692] == 43692 && 
b[43693] == 43693 && 
b[43694] == 43694 && 
b[43695] == 43695 && 
b[43696] == 43696 && 
b[43697] == 43697 && 
b[43698] == 43698 && 
b[43699] == 43699 && 
b[43700] == 43700 && 
b[43701] == 43701 && 
b[43702] == 43702 && 
b[43703] == 43703 && 
b[43704] == 43704 && 
b[43705] == 43705 && 
b[43706] == 43706 && 
b[43707] == 43707 && 
b[43708] == 43708 && 
b[43709] == 43709 && 
b[43710] == 43710 && 
b[43711] == 43711 && 
b[43712] == 43712 && 
b[43713] == 43713 && 
b[43714] == 43714 && 
b[43715] == 43715 && 
b[43716] == 43716 && 
b[43717] == 43717 && 
b[43718] == 43718 && 
b[43719] == 43719 && 
b[43720] == 43720 && 
b[43721] == 43721 && 
b[43722] == 43722 && 
b[43723] == 43723 && 
b[43724] == 43724 && 
b[43725] == 43725 && 
b[43726] == 43726 && 
b[43727] == 43727 && 
b[43728] == 43728 && 
b[43729] == 43729 && 
b[43730] == 43730 && 
b[43731] == 43731 && 
b[43732] == 43732 && 
b[43733] == 43733 && 
b[43734] == 43734 && 
b[43735] == 43735 && 
b[43736] == 43736 && 
b[43737] == 43737 && 
b[43738] == 43738 && 
b[43739] == 43739 && 
b[43740] == 43740 && 
b[43741] == 43741 && 
b[43742] == 43742 && 
b[43743] == 43743 && 
b[43744] == 43744 && 
b[43745] == 43745 && 
b[43746] == 43746 && 
b[43747] == 43747 && 
b[43748] == 43748 && 
b[43749] == 43749 && 
b[43750] == 43750 && 
b[43751] == 43751 && 
b[43752] == 43752 && 
b[43753] == 43753 && 
b[43754] == 43754 && 
b[43755] == 43755 && 
b[43756] == 43756 && 
b[43757] == 43757 && 
b[43758] == 43758 && 
b[43759] == 43759 && 
b[43760] == 43760 && 
b[43761] == 43761 && 
b[43762] == 43762 && 
b[43763] == 43763 && 
b[43764] == 43764 && 
b[43765] == 43765 && 
b[43766] == 43766 && 
b[43767] == 43767 && 
b[43768] == 43768 && 
b[43769] == 43769 && 
b[43770] == 43770 && 
b[43771] == 43771 && 
b[43772] == 43772 && 
b[43773] == 43773 && 
b[43774] == 43774 && 
b[43775] == 43775 && 
b[43776] == 43776 && 
b[43777] == 43777 && 
b[43778] == 43778 && 
b[43779] == 43779 && 
b[43780] == 43780 && 
b[43781] == 43781 && 
b[43782] == 43782 && 
b[43783] == 43783 && 
b[43784] == 43784 && 
b[43785] == 43785 && 
b[43786] == 43786 && 
b[43787] == 43787 && 
b[43788] == 43788 && 
b[43789] == 43789 && 
b[43790] == 43790 && 
b[43791] == 43791 && 
b[43792] == 43792 && 
b[43793] == 43793 && 
b[43794] == 43794 && 
b[43795] == 43795 && 
b[43796] == 43796 && 
b[43797] == 43797 && 
b[43798] == 43798 && 
b[43799] == 43799 && 
b[43800] == 43800 && 
b[43801] == 43801 && 
b[43802] == 43802 && 
b[43803] == 43803 && 
b[43804] == 43804 && 
b[43805] == 43805 && 
b[43806] == 43806 && 
b[43807] == 43807 && 
b[43808] == 43808 && 
b[43809] == 43809 && 
b[43810] == 43810 && 
b[43811] == 43811 && 
b[43812] == 43812 && 
b[43813] == 43813 && 
b[43814] == 43814 && 
b[43815] == 43815 && 
b[43816] == 43816 && 
b[43817] == 43817 && 
b[43818] == 43818 && 
b[43819] == 43819 && 
b[43820] == 43820 && 
b[43821] == 43821 && 
b[43822] == 43822 && 
b[43823] == 43823 && 
b[43824] == 43824 && 
b[43825] == 43825 && 
b[43826] == 43826 && 
b[43827] == 43827 && 
b[43828] == 43828 && 
b[43829] == 43829 && 
b[43830] == 43830 && 
b[43831] == 43831 && 
b[43832] == 43832 && 
b[43833] == 43833 && 
b[43834] == 43834 && 
b[43835] == 43835 && 
b[43836] == 43836 && 
b[43837] == 43837 && 
b[43838] == 43838 && 
b[43839] == 43839 && 
b[43840] == 43840 && 
b[43841] == 43841 && 
b[43842] == 43842 && 
b[43843] == 43843 && 
b[43844] == 43844 && 
b[43845] == 43845 && 
b[43846] == 43846 && 
b[43847] == 43847 && 
b[43848] == 43848 && 
b[43849] == 43849 && 
b[43850] == 43850 && 
b[43851] == 43851 && 
b[43852] == 43852 && 
b[43853] == 43853 && 
b[43854] == 43854 && 
b[43855] == 43855 && 
b[43856] == 43856 && 
b[43857] == 43857 && 
b[43858] == 43858 && 
b[43859] == 43859 && 
b[43860] == 43860 && 
b[43861] == 43861 && 
b[43862] == 43862 && 
b[43863] == 43863 && 
b[43864] == 43864 && 
b[43865] == 43865 && 
b[43866] == 43866 && 
b[43867] == 43867 && 
b[43868] == 43868 && 
b[43869] == 43869 && 
b[43870] == 43870 && 
b[43871] == 43871 && 
b[43872] == 43872 && 
b[43873] == 43873 && 
b[43874] == 43874 && 
b[43875] == 43875 && 
b[43876] == 43876 && 
b[43877] == 43877 && 
b[43878] == 43878 && 
b[43879] == 43879 && 
b[43880] == 43880 && 
b[43881] == 43881 && 
b[43882] == 43882 && 
b[43883] == 43883 && 
b[43884] == 43884 && 
b[43885] == 43885 && 
b[43886] == 43886 && 
b[43887] == 43887 && 
b[43888] == 43888 && 
b[43889] == 43889 && 
b[43890] == 43890 && 
b[43891] == 43891 && 
b[43892] == 43892 && 
b[43893] == 43893 && 
b[43894] == 43894 && 
b[43895] == 43895 && 
b[43896] == 43896 && 
b[43897] == 43897 && 
b[43898] == 43898 && 
b[43899] == 43899 && 
b[43900] == 43900 && 
b[43901] == 43901 && 
b[43902] == 43902 && 
b[43903] == 43903 && 
b[43904] == 43904 && 
b[43905] == 43905 && 
b[43906] == 43906 && 
b[43907] == 43907 && 
b[43908] == 43908 && 
b[43909] == 43909 && 
b[43910] == 43910 && 
b[43911] == 43911 && 
b[43912] == 43912 && 
b[43913] == 43913 && 
b[43914] == 43914 && 
b[43915] == 43915 && 
b[43916] == 43916 && 
b[43917] == 43917 && 
b[43918] == 43918 && 
b[43919] == 43919 && 
b[43920] == 43920 && 
b[43921] == 43921 && 
b[43922] == 43922 && 
b[43923] == 43923 && 
b[43924] == 43924 && 
b[43925] == 43925 && 
b[43926] == 43926 && 
b[43927] == 43927 && 
b[43928] == 43928 && 
b[43929] == 43929 && 
b[43930] == 43930 && 
b[43931] == 43931 && 
b[43932] == 43932 && 
b[43933] == 43933 && 
b[43934] == 43934 && 
b[43935] == 43935 && 
b[43936] == 43936 && 
b[43937] == 43937 && 
b[43938] == 43938 && 
b[43939] == 43939 && 
b[43940] == 43940 && 
b[43941] == 43941 && 
b[43942] == 43942 && 
b[43943] == 43943 && 
b[43944] == 43944 && 
b[43945] == 43945 && 
b[43946] == 43946 && 
b[43947] == 43947 && 
b[43948] == 43948 && 
b[43949] == 43949 && 
b[43950] == 43950 && 
b[43951] == 43951 && 
b[43952] == 43952 && 
b[43953] == 43953 && 
b[43954] == 43954 && 
b[43955] == 43955 && 
b[43956] == 43956 && 
b[43957] == 43957 && 
b[43958] == 43958 && 
b[43959] == 43959 && 
b[43960] == 43960 && 
b[43961] == 43961 && 
b[43962] == 43962 && 
b[43963] == 43963 && 
b[43964] == 43964 && 
b[43965] == 43965 && 
b[43966] == 43966 && 
b[43967] == 43967 && 
b[43968] == 43968 && 
b[43969] == 43969 && 
b[43970] == 43970 && 
b[43971] == 43971 && 
b[43972] == 43972 && 
b[43973] == 43973 && 
b[43974] == 43974 && 
b[43975] == 43975 && 
b[43976] == 43976 && 
b[43977] == 43977 && 
b[43978] == 43978 && 
b[43979] == 43979 && 
b[43980] == 43980 && 
b[43981] == 43981 && 
b[43982] == 43982 && 
b[43983] == 43983 && 
b[43984] == 43984 && 
b[43985] == 43985 && 
b[43986] == 43986 && 
b[43987] == 43987 && 
b[43988] == 43988 && 
b[43989] == 43989 && 
b[43990] == 43990 && 
b[43991] == 43991 && 
b[43992] == 43992 && 
b[43993] == 43993 && 
b[43994] == 43994 && 
b[43995] == 43995 && 
b[43996] == 43996 && 
b[43997] == 43997 && 
b[43998] == 43998 && 
b[43999] == 43999 && 
b[44000] == 44000 && 
b[44001] == 44001 && 
b[44002] == 44002 && 
b[44003] == 44003 && 
b[44004] == 44004 && 
b[44005] == 44005 && 
b[44006] == 44006 && 
b[44007] == 44007 && 
b[44008] == 44008 && 
b[44009] == 44009 && 
b[44010] == 44010 && 
b[44011] == 44011 && 
b[44012] == 44012 && 
b[44013] == 44013 && 
b[44014] == 44014 && 
b[44015] == 44015 && 
b[44016] == 44016 && 
b[44017] == 44017 && 
b[44018] == 44018 && 
b[44019] == 44019 && 
b[44020] == 44020 && 
b[44021] == 44021 && 
b[44022] == 44022 && 
b[44023] == 44023 && 
b[44024] == 44024 && 
b[44025] == 44025 && 
b[44026] == 44026 && 
b[44027] == 44027 && 
b[44028] == 44028 && 
b[44029] == 44029 && 
b[44030] == 44030 && 
b[44031] == 44031 && 
b[44032] == 44032 && 
b[44033] == 44033 && 
b[44034] == 44034 && 
b[44035] == 44035 && 
b[44036] == 44036 && 
b[44037] == 44037 && 
b[44038] == 44038 && 
b[44039] == 44039 && 
b[44040] == 44040 && 
b[44041] == 44041 && 
b[44042] == 44042 && 
b[44043] == 44043 && 
b[44044] == 44044 && 
b[44045] == 44045 && 
b[44046] == 44046 && 
b[44047] == 44047 && 
b[44048] == 44048 && 
b[44049] == 44049 && 
b[44050] == 44050 && 
b[44051] == 44051 && 
b[44052] == 44052 && 
b[44053] == 44053 && 
b[44054] == 44054 && 
b[44055] == 44055 && 
b[44056] == 44056 && 
b[44057] == 44057 && 
b[44058] == 44058 && 
b[44059] == 44059 && 
b[44060] == 44060 && 
b[44061] == 44061 && 
b[44062] == 44062 && 
b[44063] == 44063 && 
b[44064] == 44064 && 
b[44065] == 44065 && 
b[44066] == 44066 && 
b[44067] == 44067 && 
b[44068] == 44068 && 
b[44069] == 44069 && 
b[44070] == 44070 && 
b[44071] == 44071 && 
b[44072] == 44072 && 
b[44073] == 44073 && 
b[44074] == 44074 && 
b[44075] == 44075 && 
b[44076] == 44076 && 
b[44077] == 44077 && 
b[44078] == 44078 && 
b[44079] == 44079 && 
b[44080] == 44080 && 
b[44081] == 44081 && 
b[44082] == 44082 && 
b[44083] == 44083 && 
b[44084] == 44084 && 
b[44085] == 44085 && 
b[44086] == 44086 && 
b[44087] == 44087 && 
b[44088] == 44088 && 
b[44089] == 44089 && 
b[44090] == 44090 && 
b[44091] == 44091 && 
b[44092] == 44092 && 
b[44093] == 44093 && 
b[44094] == 44094 && 
b[44095] == 44095 && 
b[44096] == 44096 && 
b[44097] == 44097 && 
b[44098] == 44098 && 
b[44099] == 44099 && 
b[44100] == 44100 && 
b[44101] == 44101 && 
b[44102] == 44102 && 
b[44103] == 44103 && 
b[44104] == 44104 && 
b[44105] == 44105 && 
b[44106] == 44106 && 
b[44107] == 44107 && 
b[44108] == 44108 && 
b[44109] == 44109 && 
b[44110] == 44110 && 
b[44111] == 44111 && 
b[44112] == 44112 && 
b[44113] == 44113 && 
b[44114] == 44114 && 
b[44115] == 44115 && 
b[44116] == 44116 && 
b[44117] == 44117 && 
b[44118] == 44118 && 
b[44119] == 44119 && 
b[44120] == 44120 && 
b[44121] == 44121 && 
b[44122] == 44122 && 
b[44123] == 44123 && 
b[44124] == 44124 && 
b[44125] == 44125 && 
b[44126] == 44126 && 
b[44127] == 44127 && 
b[44128] == 44128 && 
b[44129] == 44129 && 
b[44130] == 44130 && 
b[44131] == 44131 && 
b[44132] == 44132 && 
b[44133] == 44133 && 
b[44134] == 44134 && 
b[44135] == 44135 && 
b[44136] == 44136 && 
b[44137] == 44137 && 
b[44138] == 44138 && 
b[44139] == 44139 && 
b[44140] == 44140 && 
b[44141] == 44141 && 
b[44142] == 44142 && 
b[44143] == 44143 && 
b[44144] == 44144 && 
b[44145] == 44145 && 
b[44146] == 44146 && 
b[44147] == 44147 && 
b[44148] == 44148 && 
b[44149] == 44149 && 
b[44150] == 44150 && 
b[44151] == 44151 && 
b[44152] == 44152 && 
b[44153] == 44153 && 
b[44154] == 44154 && 
b[44155] == 44155 && 
b[44156] == 44156 && 
b[44157] == 44157 && 
b[44158] == 44158 && 
b[44159] == 44159 && 
b[44160] == 44160 && 
b[44161] == 44161 && 
b[44162] == 44162 && 
b[44163] == 44163 && 
b[44164] == 44164 && 
b[44165] == 44165 && 
b[44166] == 44166 && 
b[44167] == 44167 && 
b[44168] == 44168 && 
b[44169] == 44169 && 
b[44170] == 44170 && 
b[44171] == 44171 && 
b[44172] == 44172 && 
b[44173] == 44173 && 
b[44174] == 44174 && 
b[44175] == 44175 && 
b[44176] == 44176 && 
b[44177] == 44177 && 
b[44178] == 44178 && 
b[44179] == 44179 && 
b[44180] == 44180 && 
b[44181] == 44181 && 
b[44182] == 44182 && 
b[44183] == 44183 && 
b[44184] == 44184 && 
b[44185] == 44185 && 
b[44186] == 44186 && 
b[44187] == 44187 && 
b[44188] == 44188 && 
b[44189] == 44189 && 
b[44190] == 44190 && 
b[44191] == 44191 && 
b[44192] == 44192 && 
b[44193] == 44193 && 
b[44194] == 44194 && 
b[44195] == 44195 && 
b[44196] == 44196 && 
b[44197] == 44197 && 
b[44198] == 44198 && 
b[44199] == 44199 && 
b[44200] == 44200 && 
b[44201] == 44201 && 
b[44202] == 44202 && 
b[44203] == 44203 && 
b[44204] == 44204 && 
b[44205] == 44205 && 
b[44206] == 44206 && 
b[44207] == 44207 && 
b[44208] == 44208 && 
b[44209] == 44209 && 
b[44210] == 44210 && 
b[44211] == 44211 && 
b[44212] == 44212 && 
b[44213] == 44213 && 
b[44214] == 44214 && 
b[44215] == 44215 && 
b[44216] == 44216 && 
b[44217] == 44217 && 
b[44218] == 44218 && 
b[44219] == 44219 && 
b[44220] == 44220 && 
b[44221] == 44221 && 
b[44222] == 44222 && 
b[44223] == 44223 && 
b[44224] == 44224 && 
b[44225] == 44225 && 
b[44226] == 44226 && 
b[44227] == 44227 && 
b[44228] == 44228 && 
b[44229] == 44229 && 
b[44230] == 44230 && 
b[44231] == 44231 && 
b[44232] == 44232 && 
b[44233] == 44233 && 
b[44234] == 44234 && 
b[44235] == 44235 && 
b[44236] == 44236 && 
b[44237] == 44237 && 
b[44238] == 44238 && 
b[44239] == 44239 && 
b[44240] == 44240 && 
b[44241] == 44241 && 
b[44242] == 44242 && 
b[44243] == 44243 && 
b[44244] == 44244 && 
b[44245] == 44245 && 
b[44246] == 44246 && 
b[44247] == 44247 && 
b[44248] == 44248 && 
b[44249] == 44249 && 
b[44250] == 44250 && 
b[44251] == 44251 && 
b[44252] == 44252 && 
b[44253] == 44253 && 
b[44254] == 44254 && 
b[44255] == 44255 && 
b[44256] == 44256 && 
b[44257] == 44257 && 
b[44258] == 44258 && 
b[44259] == 44259 && 
b[44260] == 44260 && 
b[44261] == 44261 && 
b[44262] == 44262 && 
b[44263] == 44263 && 
b[44264] == 44264 && 
b[44265] == 44265 && 
b[44266] == 44266 && 
b[44267] == 44267 && 
b[44268] == 44268 && 
b[44269] == 44269 && 
b[44270] == 44270 && 
b[44271] == 44271 && 
b[44272] == 44272 && 
b[44273] == 44273 && 
b[44274] == 44274 && 
b[44275] == 44275 && 
b[44276] == 44276 && 
b[44277] == 44277 && 
b[44278] == 44278 && 
b[44279] == 44279 && 
b[44280] == 44280 && 
b[44281] == 44281 && 
b[44282] == 44282 && 
b[44283] == 44283 && 
b[44284] == 44284 && 
b[44285] == 44285 && 
b[44286] == 44286 && 
b[44287] == 44287 && 
b[44288] == 44288 && 
b[44289] == 44289 && 
b[44290] == 44290 && 
b[44291] == 44291 && 
b[44292] == 44292 && 
b[44293] == 44293 && 
b[44294] == 44294 && 
b[44295] == 44295 && 
b[44296] == 44296 && 
b[44297] == 44297 && 
b[44298] == 44298 && 
b[44299] == 44299 && 
b[44300] == 44300 && 
b[44301] == 44301 && 
b[44302] == 44302 && 
b[44303] == 44303 && 
b[44304] == 44304 && 
b[44305] == 44305 && 
b[44306] == 44306 && 
b[44307] == 44307 && 
b[44308] == 44308 && 
b[44309] == 44309 && 
b[44310] == 44310 && 
b[44311] == 44311 && 
b[44312] == 44312 && 
b[44313] == 44313 && 
b[44314] == 44314 && 
b[44315] == 44315 && 
b[44316] == 44316 && 
b[44317] == 44317 && 
b[44318] == 44318 && 
b[44319] == 44319 && 
b[44320] == 44320 && 
b[44321] == 44321 && 
b[44322] == 44322 && 
b[44323] == 44323 && 
b[44324] == 44324 && 
b[44325] == 44325 && 
b[44326] == 44326 && 
b[44327] == 44327 && 
b[44328] == 44328 && 
b[44329] == 44329 && 
b[44330] == 44330 && 
b[44331] == 44331 && 
b[44332] == 44332 && 
b[44333] == 44333 && 
b[44334] == 44334 && 
b[44335] == 44335 && 
b[44336] == 44336 && 
b[44337] == 44337 && 
b[44338] == 44338 && 
b[44339] == 44339 && 
b[44340] == 44340 && 
b[44341] == 44341 && 
b[44342] == 44342 && 
b[44343] == 44343 && 
b[44344] == 44344 && 
b[44345] == 44345 && 
b[44346] == 44346 && 
b[44347] == 44347 && 
b[44348] == 44348 && 
b[44349] == 44349 && 
b[44350] == 44350 && 
b[44351] == 44351 && 
b[44352] == 44352 && 
b[44353] == 44353 && 
b[44354] == 44354 && 
b[44355] == 44355 && 
b[44356] == 44356 && 
b[44357] == 44357 && 
b[44358] == 44358 && 
b[44359] == 44359 && 
b[44360] == 44360 && 
b[44361] == 44361 && 
b[44362] == 44362 && 
b[44363] == 44363 && 
b[44364] == 44364 && 
b[44365] == 44365 && 
b[44366] == 44366 && 
b[44367] == 44367 && 
b[44368] == 44368 && 
b[44369] == 44369 && 
b[44370] == 44370 && 
b[44371] == 44371 && 
b[44372] == 44372 && 
b[44373] == 44373 && 
b[44374] == 44374 && 
b[44375] == 44375 && 
b[44376] == 44376 && 
b[44377] == 44377 && 
b[44378] == 44378 && 
b[44379] == 44379 && 
b[44380] == 44380 && 
b[44381] == 44381 && 
b[44382] == 44382 && 
b[44383] == 44383 && 
b[44384] == 44384 && 
b[44385] == 44385 && 
b[44386] == 44386 && 
b[44387] == 44387 && 
b[44388] == 44388 && 
b[44389] == 44389 && 
b[44390] == 44390 && 
b[44391] == 44391 && 
b[44392] == 44392 && 
b[44393] == 44393 && 
b[44394] == 44394 && 
b[44395] == 44395 && 
b[44396] == 44396 && 
b[44397] == 44397 && 
b[44398] == 44398 && 
b[44399] == 44399 && 
b[44400] == 44400 && 
b[44401] == 44401 && 
b[44402] == 44402 && 
b[44403] == 44403 && 
b[44404] == 44404 && 
b[44405] == 44405 && 
b[44406] == 44406 && 
b[44407] == 44407 && 
b[44408] == 44408 && 
b[44409] == 44409 && 
b[44410] == 44410 && 
b[44411] == 44411 && 
b[44412] == 44412 && 
b[44413] == 44413 && 
b[44414] == 44414 && 
b[44415] == 44415 && 
b[44416] == 44416 && 
b[44417] == 44417 && 
b[44418] == 44418 && 
b[44419] == 44419 && 
b[44420] == 44420 && 
b[44421] == 44421 && 
b[44422] == 44422 && 
b[44423] == 44423 && 
b[44424] == 44424 && 
b[44425] == 44425 && 
b[44426] == 44426 && 
b[44427] == 44427 && 
b[44428] == 44428 && 
b[44429] == 44429 && 
b[44430] == 44430 && 
b[44431] == 44431 && 
b[44432] == 44432 && 
b[44433] == 44433 && 
b[44434] == 44434 && 
b[44435] == 44435 && 
b[44436] == 44436 && 
b[44437] == 44437 && 
b[44438] == 44438 && 
b[44439] == 44439 && 
b[44440] == 44440 && 
b[44441] == 44441 && 
b[44442] == 44442 && 
b[44443] == 44443 && 
b[44444] == 44444 && 
b[44445] == 44445 && 
b[44446] == 44446 && 
b[44447] == 44447 && 
b[44448] == 44448 && 
b[44449] == 44449 && 
b[44450] == 44450 && 
b[44451] == 44451 && 
b[44452] == 44452 && 
b[44453] == 44453 && 
b[44454] == 44454 && 
b[44455] == 44455 && 
b[44456] == 44456 && 
b[44457] == 44457 && 
b[44458] == 44458 && 
b[44459] == 44459 && 
b[44460] == 44460 && 
b[44461] == 44461 && 
b[44462] == 44462 && 
b[44463] == 44463 && 
b[44464] == 44464 && 
b[44465] == 44465 && 
b[44466] == 44466 && 
b[44467] == 44467 && 
b[44468] == 44468 && 
b[44469] == 44469 && 
b[44470] == 44470 && 
b[44471] == 44471 && 
b[44472] == 44472 && 
b[44473] == 44473 && 
b[44474] == 44474 && 
b[44475] == 44475 && 
b[44476] == 44476 && 
b[44477] == 44477 && 
b[44478] == 44478 && 
b[44479] == 44479 && 
b[44480] == 44480 && 
b[44481] == 44481 && 
b[44482] == 44482 && 
b[44483] == 44483 && 
b[44484] == 44484 && 
b[44485] == 44485 && 
b[44486] == 44486 && 
b[44487] == 44487 && 
b[44488] == 44488 && 
b[44489] == 44489 && 
b[44490] == 44490 && 
b[44491] == 44491 && 
b[44492] == 44492 && 
b[44493] == 44493 && 
b[44494] == 44494 && 
b[44495] == 44495 && 
b[44496] == 44496 && 
b[44497] == 44497 && 
b[44498] == 44498 && 
b[44499] == 44499 && 
b[44500] == 44500 && 
b[44501] == 44501 && 
b[44502] == 44502 && 
b[44503] == 44503 && 
b[44504] == 44504 && 
b[44505] == 44505 && 
b[44506] == 44506 && 
b[44507] == 44507 && 
b[44508] == 44508 && 
b[44509] == 44509 && 
b[44510] == 44510 && 
b[44511] == 44511 && 
b[44512] == 44512 && 
b[44513] == 44513 && 
b[44514] == 44514 && 
b[44515] == 44515 && 
b[44516] == 44516 && 
b[44517] == 44517 && 
b[44518] == 44518 && 
b[44519] == 44519 && 
b[44520] == 44520 && 
b[44521] == 44521 && 
b[44522] == 44522 && 
b[44523] == 44523 && 
b[44524] == 44524 && 
b[44525] == 44525 && 
b[44526] == 44526 && 
b[44527] == 44527 && 
b[44528] == 44528 && 
b[44529] == 44529 && 
b[44530] == 44530 && 
b[44531] == 44531 && 
b[44532] == 44532 && 
b[44533] == 44533 && 
b[44534] == 44534 && 
b[44535] == 44535 && 
b[44536] == 44536 && 
b[44537] == 44537 && 
b[44538] == 44538 && 
b[44539] == 44539 && 
b[44540] == 44540 && 
b[44541] == 44541 && 
b[44542] == 44542 && 
b[44543] == 44543 && 
b[44544] == 44544 && 
b[44545] == 44545 && 
b[44546] == 44546 && 
b[44547] == 44547 && 
b[44548] == 44548 && 
b[44549] == 44549 && 
b[44550] == 44550 && 
b[44551] == 44551 && 
b[44552] == 44552 && 
b[44553] == 44553 && 
b[44554] == 44554 && 
b[44555] == 44555 && 
b[44556] == 44556 && 
b[44557] == 44557 && 
b[44558] == 44558 && 
b[44559] == 44559 && 
b[44560] == 44560 && 
b[44561] == 44561 && 
b[44562] == 44562 && 
b[44563] == 44563 && 
b[44564] == 44564 && 
b[44565] == 44565 && 
b[44566] == 44566 && 
b[44567] == 44567 && 
b[44568] == 44568 && 
b[44569] == 44569 && 
b[44570] == 44570 && 
b[44571] == 44571 && 
b[44572] == 44572 && 
b[44573] == 44573 && 
b[44574] == 44574 && 
b[44575] == 44575 && 
b[44576] == 44576 && 
b[44577] == 44577 && 
b[44578] == 44578 && 
b[44579] == 44579 && 
b[44580] == 44580 && 
b[44581] == 44581 && 
b[44582] == 44582 && 
b[44583] == 44583 && 
b[44584] == 44584 && 
b[44585] == 44585 && 
b[44586] == 44586 && 
b[44587] == 44587 && 
b[44588] == 44588 && 
b[44589] == 44589 && 
b[44590] == 44590 && 
b[44591] == 44591 && 
b[44592] == 44592 && 
b[44593] == 44593 && 
b[44594] == 44594 && 
b[44595] == 44595 && 
b[44596] == 44596 && 
b[44597] == 44597 && 
b[44598] == 44598 && 
b[44599] == 44599 && 
b[44600] == 44600 && 
b[44601] == 44601 && 
b[44602] == 44602 && 
b[44603] == 44603 && 
b[44604] == 44604 && 
b[44605] == 44605 && 
b[44606] == 44606 && 
b[44607] == 44607 && 
b[44608] == 44608 && 
b[44609] == 44609 && 
b[44610] == 44610 && 
b[44611] == 44611 && 
b[44612] == 44612 && 
b[44613] == 44613 && 
b[44614] == 44614 && 
b[44615] == 44615 && 
b[44616] == 44616 && 
b[44617] == 44617 && 
b[44618] == 44618 && 
b[44619] == 44619 && 
b[44620] == 44620 && 
b[44621] == 44621 && 
b[44622] == 44622 && 
b[44623] == 44623 && 
b[44624] == 44624 && 
b[44625] == 44625 && 
b[44626] == 44626 && 
b[44627] == 44627 && 
b[44628] == 44628 && 
b[44629] == 44629 && 
b[44630] == 44630 && 
b[44631] == 44631 && 
b[44632] == 44632 && 
b[44633] == 44633 && 
b[44634] == 44634 && 
b[44635] == 44635 && 
b[44636] == 44636 && 
b[44637] == 44637 && 
b[44638] == 44638 && 
b[44639] == 44639 && 
b[44640] == 44640 && 
b[44641] == 44641 && 
b[44642] == 44642 && 
b[44643] == 44643 && 
b[44644] == 44644 && 
b[44645] == 44645 && 
b[44646] == 44646 && 
b[44647] == 44647 && 
b[44648] == 44648 && 
b[44649] == 44649 && 
b[44650] == 44650 && 
b[44651] == 44651 && 
b[44652] == 44652 && 
b[44653] == 44653 && 
b[44654] == 44654 && 
b[44655] == 44655 && 
b[44656] == 44656 && 
b[44657] == 44657 && 
b[44658] == 44658 && 
b[44659] == 44659 && 
b[44660] == 44660 && 
b[44661] == 44661 && 
b[44662] == 44662 && 
b[44663] == 44663 && 
b[44664] == 44664 && 
b[44665] == 44665 && 
b[44666] == 44666 && 
b[44667] == 44667 && 
b[44668] == 44668 && 
b[44669] == 44669 && 
b[44670] == 44670 && 
b[44671] == 44671 && 
b[44672] == 44672 && 
b[44673] == 44673 && 
b[44674] == 44674 && 
b[44675] == 44675 && 
b[44676] == 44676 && 
b[44677] == 44677 && 
b[44678] == 44678 && 
b[44679] == 44679 && 
b[44680] == 44680 && 
b[44681] == 44681 && 
b[44682] == 44682 && 
b[44683] == 44683 && 
b[44684] == 44684 && 
b[44685] == 44685 && 
b[44686] == 44686 && 
b[44687] == 44687 && 
b[44688] == 44688 && 
b[44689] == 44689 && 
b[44690] == 44690 && 
b[44691] == 44691 && 
b[44692] == 44692 && 
b[44693] == 44693 && 
b[44694] == 44694 && 
b[44695] == 44695 && 
b[44696] == 44696 && 
b[44697] == 44697 && 
b[44698] == 44698 && 
b[44699] == 44699 && 
b[44700] == 44700 && 
b[44701] == 44701 && 
b[44702] == 44702 && 
b[44703] == 44703 && 
b[44704] == 44704 && 
b[44705] == 44705 && 
b[44706] == 44706 && 
b[44707] == 44707 && 
b[44708] == 44708 && 
b[44709] == 44709 && 
b[44710] == 44710 && 
b[44711] == 44711 && 
b[44712] == 44712 && 
b[44713] == 44713 && 
b[44714] == 44714 && 
b[44715] == 44715 && 
b[44716] == 44716 && 
b[44717] == 44717 && 
b[44718] == 44718 && 
b[44719] == 44719 && 
b[44720] == 44720 && 
b[44721] == 44721 && 
b[44722] == 44722 && 
b[44723] == 44723 && 
b[44724] == 44724 && 
b[44725] == 44725 && 
b[44726] == 44726 && 
b[44727] == 44727 && 
b[44728] == 44728 && 
b[44729] == 44729 && 
b[44730] == 44730 && 
b[44731] == 44731 && 
b[44732] == 44732 && 
b[44733] == 44733 && 
b[44734] == 44734 && 
b[44735] == 44735 && 
b[44736] == 44736 && 
b[44737] == 44737 && 
b[44738] == 44738 && 
b[44739] == 44739 && 
b[44740] == 44740 && 
b[44741] == 44741 && 
b[44742] == 44742 && 
b[44743] == 44743 && 
b[44744] == 44744 && 
b[44745] == 44745 && 
b[44746] == 44746 && 
b[44747] == 44747 && 
b[44748] == 44748 && 
b[44749] == 44749 && 
b[44750] == 44750 && 
b[44751] == 44751 && 
b[44752] == 44752 && 
b[44753] == 44753 && 
b[44754] == 44754 && 
b[44755] == 44755 && 
b[44756] == 44756 && 
b[44757] == 44757 && 
b[44758] == 44758 && 
b[44759] == 44759 && 
b[44760] == 44760 && 
b[44761] == 44761 && 
b[44762] == 44762 && 
b[44763] == 44763 && 
b[44764] == 44764 && 
b[44765] == 44765 && 
b[44766] == 44766 && 
b[44767] == 44767 && 
b[44768] == 44768 && 
b[44769] == 44769 && 
b[44770] == 44770 && 
b[44771] == 44771 && 
b[44772] == 44772 && 
b[44773] == 44773 && 
b[44774] == 44774 && 
b[44775] == 44775 && 
b[44776] == 44776 && 
b[44777] == 44777 && 
b[44778] == 44778 && 
b[44779] == 44779 && 
b[44780] == 44780 && 
b[44781] == 44781 && 
b[44782] == 44782 && 
b[44783] == 44783 && 
b[44784] == 44784 && 
b[44785] == 44785 && 
b[44786] == 44786 && 
b[44787] == 44787 && 
b[44788] == 44788 && 
b[44789] == 44789 && 
b[44790] == 44790 && 
b[44791] == 44791 && 
b[44792] == 44792 && 
b[44793] == 44793 && 
b[44794] == 44794 && 
b[44795] == 44795 && 
b[44796] == 44796 && 
b[44797] == 44797 && 
b[44798] == 44798 && 
b[44799] == 44799 && 
b[44800] == 44800 && 
b[44801] == 44801 && 
b[44802] == 44802 && 
b[44803] == 44803 && 
b[44804] == 44804 && 
b[44805] == 44805 && 
b[44806] == 44806 && 
b[44807] == 44807 && 
b[44808] == 44808 && 
b[44809] == 44809 && 
b[44810] == 44810 && 
b[44811] == 44811 && 
b[44812] == 44812 && 
b[44813] == 44813 && 
b[44814] == 44814 && 
b[44815] == 44815 && 
b[44816] == 44816 && 
b[44817] == 44817 && 
b[44818] == 44818 && 
b[44819] == 44819 && 
b[44820] == 44820 && 
b[44821] == 44821 && 
b[44822] == 44822 && 
b[44823] == 44823 && 
b[44824] == 44824 && 
b[44825] == 44825 && 
b[44826] == 44826 && 
b[44827] == 44827 && 
b[44828] == 44828 && 
b[44829] == 44829 && 
b[44830] == 44830 && 
b[44831] == 44831 && 
b[44832] == 44832 && 
b[44833] == 44833 && 
b[44834] == 44834 && 
b[44835] == 44835 && 
b[44836] == 44836 && 
b[44837] == 44837 && 
b[44838] == 44838 && 
b[44839] == 44839 && 
b[44840] == 44840 && 
b[44841] == 44841 && 
b[44842] == 44842 && 
b[44843] == 44843 && 
b[44844] == 44844 && 
b[44845] == 44845 && 
b[44846] == 44846 && 
b[44847] == 44847 && 
b[44848] == 44848 && 
b[44849] == 44849 && 
b[44850] == 44850 && 
b[44851] == 44851 && 
b[44852] == 44852 && 
b[44853] == 44853 && 
b[44854] == 44854 && 
b[44855] == 44855 && 
b[44856] == 44856 && 
b[44857] == 44857 && 
b[44858] == 44858 && 
b[44859] == 44859 && 
b[44860] == 44860 && 
b[44861] == 44861 && 
b[44862] == 44862 && 
b[44863] == 44863 && 
b[44864] == 44864 && 
b[44865] == 44865 && 
b[44866] == 44866 && 
b[44867] == 44867 && 
b[44868] == 44868 && 
b[44869] == 44869 && 
b[44870] == 44870 && 
b[44871] == 44871 && 
b[44872] == 44872 && 
b[44873] == 44873 && 
b[44874] == 44874 && 
b[44875] == 44875 && 
b[44876] == 44876 && 
b[44877] == 44877 && 
b[44878] == 44878 && 
b[44879] == 44879 && 
b[44880] == 44880 && 
b[44881] == 44881 && 
b[44882] == 44882 && 
b[44883] == 44883 && 
b[44884] == 44884 && 
b[44885] == 44885 && 
b[44886] == 44886 && 
b[44887] == 44887 && 
b[44888] == 44888 && 
b[44889] == 44889 && 
b[44890] == 44890 && 
b[44891] == 44891 && 
b[44892] == 44892 && 
b[44893] == 44893 && 
b[44894] == 44894 && 
b[44895] == 44895 && 
b[44896] == 44896 && 
b[44897] == 44897 && 
b[44898] == 44898 && 
b[44899] == 44899 && 
b[44900] == 44900 && 
b[44901] == 44901 && 
b[44902] == 44902 && 
b[44903] == 44903 && 
b[44904] == 44904 && 
b[44905] == 44905 && 
b[44906] == 44906 && 
b[44907] == 44907 && 
b[44908] == 44908 && 
b[44909] == 44909 && 
b[44910] == 44910 && 
b[44911] == 44911 && 
b[44912] == 44912 && 
b[44913] == 44913 && 
b[44914] == 44914 && 
b[44915] == 44915 && 
b[44916] == 44916 && 
b[44917] == 44917 && 
b[44918] == 44918 && 
b[44919] == 44919 && 
b[44920] == 44920 && 
b[44921] == 44921 && 
b[44922] == 44922 && 
b[44923] == 44923 && 
b[44924] == 44924 && 
b[44925] == 44925 && 
b[44926] == 44926 && 
b[44927] == 44927 && 
b[44928] == 44928 && 
b[44929] == 44929 && 
b[44930] == 44930 && 
b[44931] == 44931 && 
b[44932] == 44932 && 
b[44933] == 44933 && 
b[44934] == 44934 && 
b[44935] == 44935 && 
b[44936] == 44936 && 
b[44937] == 44937 && 
b[44938] == 44938 && 
b[44939] == 44939 && 
b[44940] == 44940 && 
b[44941] == 44941 && 
b[44942] == 44942 && 
b[44943] == 44943 && 
b[44944] == 44944 && 
b[44945] == 44945 && 
b[44946] == 44946 && 
b[44947] == 44947 && 
b[44948] == 44948 && 
b[44949] == 44949 && 
b[44950] == 44950 && 
b[44951] == 44951 && 
b[44952] == 44952 && 
b[44953] == 44953 && 
b[44954] == 44954 && 
b[44955] == 44955 && 
b[44956] == 44956 && 
b[44957] == 44957 && 
b[44958] == 44958 && 
b[44959] == 44959 && 
b[44960] == 44960 && 
b[44961] == 44961 && 
b[44962] == 44962 && 
b[44963] == 44963 && 
b[44964] == 44964 && 
b[44965] == 44965 && 
b[44966] == 44966 && 
b[44967] == 44967 && 
b[44968] == 44968 && 
b[44969] == 44969 && 
b[44970] == 44970 && 
b[44971] == 44971 && 
b[44972] == 44972 && 
b[44973] == 44973 && 
b[44974] == 44974 && 
b[44975] == 44975 && 
b[44976] == 44976 && 
b[44977] == 44977 && 
b[44978] == 44978 && 
b[44979] == 44979 && 
b[44980] == 44980 && 
b[44981] == 44981 && 
b[44982] == 44982 && 
b[44983] == 44983 && 
b[44984] == 44984 && 
b[44985] == 44985 && 
b[44986] == 44986 && 
b[44987] == 44987 && 
b[44988] == 44988 && 
b[44989] == 44989 && 
b[44990] == 44990 && 
b[44991] == 44991 && 
b[44992] == 44992 && 
b[44993] == 44993 && 
b[44994] == 44994 && 
b[44995] == 44995 && 
b[44996] == 44996 && 
b[44997] == 44997 && 
b[44998] == 44998 && 
b[44999] == 44999 && 
b[45000] == 45000 && 
b[45001] == 45001 && 
b[45002] == 45002 && 
b[45003] == 45003 && 
b[45004] == 45004 && 
b[45005] == 45005 && 
b[45006] == 45006 && 
b[45007] == 45007 && 
b[45008] == 45008 && 
b[45009] == 45009 && 
b[45010] == 45010 && 
b[45011] == 45011 && 
b[45012] == 45012 && 
b[45013] == 45013 && 
b[45014] == 45014 && 
b[45015] == 45015 && 
b[45016] == 45016 && 
b[45017] == 45017 && 
b[45018] == 45018 && 
b[45019] == 45019 && 
b[45020] == 45020 && 
b[45021] == 45021 && 
b[45022] == 45022 && 
b[45023] == 45023 && 
b[45024] == 45024 && 
b[45025] == 45025 && 
b[45026] == 45026 && 
b[45027] == 45027 && 
b[45028] == 45028 && 
b[45029] == 45029 && 
b[45030] == 45030 && 
b[45031] == 45031 && 
b[45032] == 45032 && 
b[45033] == 45033 && 
b[45034] == 45034 && 
b[45035] == 45035 && 
b[45036] == 45036 && 
b[45037] == 45037 && 
b[45038] == 45038 && 
b[45039] == 45039 && 
b[45040] == 45040 && 
b[45041] == 45041 && 
b[45042] == 45042 && 
b[45043] == 45043 && 
b[45044] == 45044 && 
b[45045] == 45045 && 
b[45046] == 45046 && 
b[45047] == 45047 && 
b[45048] == 45048 && 
b[45049] == 45049 && 
b[45050] == 45050 && 
b[45051] == 45051 && 
b[45052] == 45052 && 
b[45053] == 45053 && 
b[45054] == 45054 && 
b[45055] == 45055 && 
b[45056] == 45056 && 
b[45057] == 45057 && 
b[45058] == 45058 && 
b[45059] == 45059 && 
b[45060] == 45060 && 
b[45061] == 45061 && 
b[45062] == 45062 && 
b[45063] == 45063 && 
b[45064] == 45064 && 
b[45065] == 45065 && 
b[45066] == 45066 && 
b[45067] == 45067 && 
b[45068] == 45068 && 
b[45069] == 45069 && 
b[45070] == 45070 && 
b[45071] == 45071 && 
b[45072] == 45072 && 
b[45073] == 45073 && 
b[45074] == 45074 && 
b[45075] == 45075 && 
b[45076] == 45076 && 
b[45077] == 45077 && 
b[45078] == 45078 && 
b[45079] == 45079 && 
b[45080] == 45080 && 
b[45081] == 45081 && 
b[45082] == 45082 && 
b[45083] == 45083 && 
b[45084] == 45084 && 
b[45085] == 45085 && 
b[45086] == 45086 && 
b[45087] == 45087 && 
b[45088] == 45088 && 
b[45089] == 45089 && 
b[45090] == 45090 && 
b[45091] == 45091 && 
b[45092] == 45092 && 
b[45093] == 45093 && 
b[45094] == 45094 && 
b[45095] == 45095 && 
b[45096] == 45096 && 
b[45097] == 45097 && 
b[45098] == 45098 && 
b[45099] == 45099 && 
b[45100] == 45100 && 
b[45101] == 45101 && 
b[45102] == 45102 && 
b[45103] == 45103 && 
b[45104] == 45104 && 
b[45105] == 45105 && 
b[45106] == 45106 && 
b[45107] == 45107 && 
b[45108] == 45108 && 
b[45109] == 45109 && 
b[45110] == 45110 && 
b[45111] == 45111 && 
b[45112] == 45112 && 
b[45113] == 45113 && 
b[45114] == 45114 && 
b[45115] == 45115 && 
b[45116] == 45116 && 
b[45117] == 45117 && 
b[45118] == 45118 && 
b[45119] == 45119 && 
b[45120] == 45120 && 
b[45121] == 45121 && 
b[45122] == 45122 && 
b[45123] == 45123 && 
b[45124] == 45124 && 
b[45125] == 45125 && 
b[45126] == 45126 && 
b[45127] == 45127 && 
b[45128] == 45128 && 
b[45129] == 45129 && 
b[45130] == 45130 && 
b[45131] == 45131 && 
b[45132] == 45132 && 
b[45133] == 45133 && 
b[45134] == 45134 && 
b[45135] == 45135 && 
b[45136] == 45136 && 
b[45137] == 45137 && 
b[45138] == 45138 && 
b[45139] == 45139 && 
b[45140] == 45140 && 
b[45141] == 45141 && 
b[45142] == 45142 && 
b[45143] == 45143 && 
b[45144] == 45144 && 
b[45145] == 45145 && 
b[45146] == 45146 && 
b[45147] == 45147 && 
b[45148] == 45148 && 
b[45149] == 45149 && 
b[45150] == 45150 && 
b[45151] == 45151 && 
b[45152] == 45152 && 
b[45153] == 45153 && 
b[45154] == 45154 && 
b[45155] == 45155 && 
b[45156] == 45156 && 
b[45157] == 45157 && 
b[45158] == 45158 && 
b[45159] == 45159 && 
b[45160] == 45160 && 
b[45161] == 45161 && 
b[45162] == 45162 && 
b[45163] == 45163 && 
b[45164] == 45164 && 
b[45165] == 45165 && 
b[45166] == 45166 && 
b[45167] == 45167 && 
b[45168] == 45168 && 
b[45169] == 45169 && 
b[45170] == 45170 && 
b[45171] == 45171 && 
b[45172] == 45172 && 
b[45173] == 45173 && 
b[45174] == 45174 && 
b[45175] == 45175 && 
b[45176] == 45176 && 
b[45177] == 45177 && 
b[45178] == 45178 && 
b[45179] == 45179 && 
b[45180] == 45180 && 
b[45181] == 45181 && 
b[45182] == 45182 && 
b[45183] == 45183 && 
b[45184] == 45184 && 
b[45185] == 45185 && 
b[45186] == 45186 && 
b[45187] == 45187 && 
b[45188] == 45188 && 
b[45189] == 45189 && 
b[45190] == 45190 && 
b[45191] == 45191 && 
b[45192] == 45192 && 
b[45193] == 45193 && 
b[45194] == 45194 && 
b[45195] == 45195 && 
b[45196] == 45196 && 
b[45197] == 45197 && 
b[45198] == 45198 && 
b[45199] == 45199 && 
b[45200] == 45200 && 
b[45201] == 45201 && 
b[45202] == 45202 && 
b[45203] == 45203 && 
b[45204] == 45204 && 
b[45205] == 45205 && 
b[45206] == 45206 && 
b[45207] == 45207 && 
b[45208] == 45208 && 
b[45209] == 45209 && 
b[45210] == 45210 && 
b[45211] == 45211 && 
b[45212] == 45212 && 
b[45213] == 45213 && 
b[45214] == 45214 && 
b[45215] == 45215 && 
b[45216] == 45216 && 
b[45217] == 45217 && 
b[45218] == 45218 && 
b[45219] == 45219 && 
b[45220] == 45220 && 
b[45221] == 45221 && 
b[45222] == 45222 && 
b[45223] == 45223 && 
b[45224] == 45224 && 
b[45225] == 45225 && 
b[45226] == 45226 && 
b[45227] == 45227 && 
b[45228] == 45228 && 
b[45229] == 45229 && 
b[45230] == 45230 && 
b[45231] == 45231 && 
b[45232] == 45232 && 
b[45233] == 45233 && 
b[45234] == 45234 && 
b[45235] == 45235 && 
b[45236] == 45236 && 
b[45237] == 45237 && 
b[45238] == 45238 && 
b[45239] == 45239 && 
b[45240] == 45240 && 
b[45241] == 45241 && 
b[45242] == 45242 && 
b[45243] == 45243 && 
b[45244] == 45244 && 
b[45245] == 45245 && 
b[45246] == 45246 && 
b[45247] == 45247 && 
b[45248] == 45248 && 
b[45249] == 45249 && 
b[45250] == 45250 && 
b[45251] == 45251 && 
b[45252] == 45252 && 
b[45253] == 45253 && 
b[45254] == 45254 && 
b[45255] == 45255 && 
b[45256] == 45256 && 
b[45257] == 45257 && 
b[45258] == 45258 && 
b[45259] == 45259 && 
b[45260] == 45260 && 
b[45261] == 45261 && 
b[45262] == 45262 && 
b[45263] == 45263 && 
b[45264] == 45264 && 
b[45265] == 45265 && 
b[45266] == 45266 && 
b[45267] == 45267 && 
b[45268] == 45268 && 
b[45269] == 45269 && 
b[45270] == 45270 && 
b[45271] == 45271 && 
b[45272] == 45272 && 
b[45273] == 45273 && 
b[45274] == 45274 && 
b[45275] == 45275 && 
b[45276] == 45276 && 
b[45277] == 45277 && 
b[45278] == 45278 && 
b[45279] == 45279 && 
b[45280] == 45280 && 
b[45281] == 45281 && 
b[45282] == 45282 && 
b[45283] == 45283 && 
b[45284] == 45284 && 
b[45285] == 45285 && 
b[45286] == 45286 && 
b[45287] == 45287 && 
b[45288] == 45288 && 
b[45289] == 45289 && 
b[45290] == 45290 && 
b[45291] == 45291 && 
b[45292] == 45292 && 
b[45293] == 45293 && 
b[45294] == 45294 && 
b[45295] == 45295 && 
b[45296] == 45296 && 
b[45297] == 45297 && 
b[45298] == 45298 && 
b[45299] == 45299 && 
b[45300] == 45300 && 
b[45301] == 45301 && 
b[45302] == 45302 && 
b[45303] == 45303 && 
b[45304] == 45304 && 
b[45305] == 45305 && 
b[45306] == 45306 && 
b[45307] == 45307 && 
b[45308] == 45308 && 
b[45309] == 45309 && 
b[45310] == 45310 && 
b[45311] == 45311 && 
b[45312] == 45312 && 
b[45313] == 45313 && 
b[45314] == 45314 && 
b[45315] == 45315 && 
b[45316] == 45316 && 
b[45317] == 45317 && 
b[45318] == 45318 && 
b[45319] == 45319 && 
b[45320] == 45320 && 
b[45321] == 45321 && 
b[45322] == 45322 && 
b[45323] == 45323 && 
b[45324] == 45324 && 
b[45325] == 45325 && 
b[45326] == 45326 && 
b[45327] == 45327 && 
b[45328] == 45328 && 
b[45329] == 45329 && 
b[45330] == 45330 && 
b[45331] == 45331 && 
b[45332] == 45332 && 
b[45333] == 45333 && 
b[45334] == 45334 && 
b[45335] == 45335 && 
b[45336] == 45336 && 
b[45337] == 45337 && 
b[45338] == 45338 && 
b[45339] == 45339 && 
b[45340] == 45340 && 
b[45341] == 45341 && 
b[45342] == 45342 && 
b[45343] == 45343 && 
b[45344] == 45344 && 
b[45345] == 45345 && 
b[45346] == 45346 && 
b[45347] == 45347 && 
b[45348] == 45348 && 
b[45349] == 45349 && 
b[45350] == 45350 && 
b[45351] == 45351 && 
b[45352] == 45352 && 
b[45353] == 45353 && 
b[45354] == 45354 && 
b[45355] == 45355 && 
b[45356] == 45356 && 
b[45357] == 45357 && 
b[45358] == 45358 && 
b[45359] == 45359 && 
b[45360] == 45360 && 
b[45361] == 45361 && 
b[45362] == 45362 && 
b[45363] == 45363 && 
b[45364] == 45364 && 
b[45365] == 45365 && 
b[45366] == 45366 && 
b[45367] == 45367 && 
b[45368] == 45368 && 
b[45369] == 45369 && 
b[45370] == 45370 && 
b[45371] == 45371 && 
b[45372] == 45372 && 
b[45373] == 45373 && 
b[45374] == 45374 && 
b[45375] == 45375 && 
b[45376] == 45376 && 
b[45377] == 45377 && 
b[45378] == 45378 && 
b[45379] == 45379 && 
b[45380] == 45380 && 
b[45381] == 45381 && 
b[45382] == 45382 && 
b[45383] == 45383 && 
b[45384] == 45384 && 
b[45385] == 45385 && 
b[45386] == 45386 && 
b[45387] == 45387 && 
b[45388] == 45388 && 
b[45389] == 45389 && 
b[45390] == 45390 && 
b[45391] == 45391 && 
b[45392] == 45392 && 
b[45393] == 45393 && 
b[45394] == 45394 && 
b[45395] == 45395 && 
b[45396] == 45396 && 
b[45397] == 45397 && 
b[45398] == 45398 && 
b[45399] == 45399 && 
b[45400] == 45400 && 
b[45401] == 45401 && 
b[45402] == 45402 && 
b[45403] == 45403 && 
b[45404] == 45404 && 
b[45405] == 45405 && 
b[45406] == 45406 && 
b[45407] == 45407 && 
b[45408] == 45408 && 
b[45409] == 45409 && 
b[45410] == 45410 && 
b[45411] == 45411 && 
b[45412] == 45412 && 
b[45413] == 45413 && 
b[45414] == 45414 && 
b[45415] == 45415 && 
b[45416] == 45416 && 
b[45417] == 45417 && 
b[45418] == 45418 && 
b[45419] == 45419 && 
b[45420] == 45420 && 
b[45421] == 45421 && 
b[45422] == 45422 && 
b[45423] == 45423 && 
b[45424] == 45424 && 
b[45425] == 45425 && 
b[45426] == 45426 && 
b[45427] == 45427 && 
b[45428] == 45428 && 
b[45429] == 45429 && 
b[45430] == 45430 && 
b[45431] == 45431 && 
b[45432] == 45432 && 
b[45433] == 45433 && 
b[45434] == 45434 && 
b[45435] == 45435 && 
b[45436] == 45436 && 
b[45437] == 45437 && 
b[45438] == 45438 && 
b[45439] == 45439 && 
b[45440] == 45440 && 
b[45441] == 45441 && 
b[45442] == 45442 && 
b[45443] == 45443 && 
b[45444] == 45444 && 
b[45445] == 45445 && 
b[45446] == 45446 && 
b[45447] == 45447 && 
b[45448] == 45448 && 
b[45449] == 45449 && 
b[45450] == 45450 && 
b[45451] == 45451 && 
b[45452] == 45452 && 
b[45453] == 45453 && 
b[45454] == 45454 && 
b[45455] == 45455 && 
b[45456] == 45456 && 
b[45457] == 45457 && 
b[45458] == 45458 && 
b[45459] == 45459 && 
b[45460] == 45460 && 
b[45461] == 45461 && 
b[45462] == 45462 && 
b[45463] == 45463 && 
b[45464] == 45464 && 
b[45465] == 45465 && 
b[45466] == 45466 && 
b[45467] == 45467 && 
b[45468] == 45468 && 
b[45469] == 45469 && 
b[45470] == 45470 && 
b[45471] == 45471 && 
b[45472] == 45472 && 
b[45473] == 45473 && 
b[45474] == 45474 && 
b[45475] == 45475 && 
b[45476] == 45476 && 
b[45477] == 45477 && 
b[45478] == 45478 && 
b[45479] == 45479 && 
b[45480] == 45480 && 
b[45481] == 45481 && 
b[45482] == 45482 && 
b[45483] == 45483 && 
b[45484] == 45484 && 
b[45485] == 45485 && 
b[45486] == 45486 && 
b[45487] == 45487 && 
b[45488] == 45488 && 
b[45489] == 45489 && 
b[45490] == 45490 && 
b[45491] == 45491 && 
b[45492] == 45492 && 
b[45493] == 45493 && 
b[45494] == 45494 && 
b[45495] == 45495 && 
b[45496] == 45496 && 
b[45497] == 45497 && 
b[45498] == 45498 && 
b[45499] == 45499 && 
b[45500] == 45500 && 
b[45501] == 45501 && 
b[45502] == 45502 && 
b[45503] == 45503 && 
b[45504] == 45504 && 
b[45505] == 45505 && 
b[45506] == 45506 && 
b[45507] == 45507 && 
b[45508] == 45508 && 
b[45509] == 45509 && 
b[45510] == 45510 && 
b[45511] == 45511 && 
b[45512] == 45512 && 
b[45513] == 45513 && 
b[45514] == 45514 && 
b[45515] == 45515 && 
b[45516] == 45516 && 
b[45517] == 45517 && 
b[45518] == 45518 && 
b[45519] == 45519 && 
b[45520] == 45520 && 
b[45521] == 45521 && 
b[45522] == 45522 && 
b[45523] == 45523 && 
b[45524] == 45524 && 
b[45525] == 45525 && 
b[45526] == 45526 && 
b[45527] == 45527 && 
b[45528] == 45528 && 
b[45529] == 45529 && 
b[45530] == 45530 && 
b[45531] == 45531 && 
b[45532] == 45532 && 
b[45533] == 45533 && 
b[45534] == 45534 && 
b[45535] == 45535 && 
b[45536] == 45536 && 
b[45537] == 45537 && 
b[45538] == 45538 && 
b[45539] == 45539 && 
b[45540] == 45540 && 
b[45541] == 45541 && 
b[45542] == 45542 && 
b[45543] == 45543 && 
b[45544] == 45544 && 
b[45545] == 45545 && 
b[45546] == 45546 && 
b[45547] == 45547 && 
b[45548] == 45548 && 
b[45549] == 45549 && 
b[45550] == 45550 && 
b[45551] == 45551 && 
b[45552] == 45552 && 
b[45553] == 45553 && 
b[45554] == 45554 && 
b[45555] == 45555 && 
b[45556] == 45556 && 
b[45557] == 45557 && 
b[45558] == 45558 && 
b[45559] == 45559 && 
b[45560] == 45560 && 
b[45561] == 45561 && 
b[45562] == 45562 && 
b[45563] == 45563 && 
b[45564] == 45564 && 
b[45565] == 45565 && 
b[45566] == 45566 && 
b[45567] == 45567 && 
b[45568] == 45568 && 
b[45569] == 45569 && 
b[45570] == 45570 && 
b[45571] == 45571 && 
b[45572] == 45572 && 
b[45573] == 45573 && 
b[45574] == 45574 && 
b[45575] == 45575 && 
b[45576] == 45576 && 
b[45577] == 45577 && 
b[45578] == 45578 && 
b[45579] == 45579 && 
b[45580] == 45580 && 
b[45581] == 45581 && 
b[45582] == 45582 && 
b[45583] == 45583 && 
b[45584] == 45584 && 
b[45585] == 45585 && 
b[45586] == 45586 && 
b[45587] == 45587 && 
b[45588] == 45588 && 
b[45589] == 45589 && 
b[45590] == 45590 && 
b[45591] == 45591 && 
b[45592] == 45592 && 
b[45593] == 45593 && 
b[45594] == 45594 && 
b[45595] == 45595 && 
b[45596] == 45596 && 
b[45597] == 45597 && 
b[45598] == 45598 && 
b[45599] == 45599 && 
b[45600] == 45600 && 
b[45601] == 45601 && 
b[45602] == 45602 && 
b[45603] == 45603 && 
b[45604] == 45604 && 
b[45605] == 45605 && 
b[45606] == 45606 && 
b[45607] == 45607 && 
b[45608] == 45608 && 
b[45609] == 45609 && 
b[45610] == 45610 && 
b[45611] == 45611 && 
b[45612] == 45612 && 
b[45613] == 45613 && 
b[45614] == 45614 && 
b[45615] == 45615 && 
b[45616] == 45616 && 
b[45617] == 45617 && 
b[45618] == 45618 && 
b[45619] == 45619 && 
b[45620] == 45620 && 
b[45621] == 45621 && 
b[45622] == 45622 && 
b[45623] == 45623 && 
b[45624] == 45624 && 
b[45625] == 45625 && 
b[45626] == 45626 && 
b[45627] == 45627 && 
b[45628] == 45628 && 
b[45629] == 45629 && 
b[45630] == 45630 && 
b[45631] == 45631 && 
b[45632] == 45632 && 
b[45633] == 45633 && 
b[45634] == 45634 && 
b[45635] == 45635 && 
b[45636] == 45636 && 
b[45637] == 45637 && 
b[45638] == 45638 && 
b[45639] == 45639 && 
b[45640] == 45640 && 
b[45641] == 45641 && 
b[45642] == 45642 && 
b[45643] == 45643 && 
b[45644] == 45644 && 
b[45645] == 45645 && 
b[45646] == 45646 && 
b[45647] == 45647 && 
b[45648] == 45648 && 
b[45649] == 45649 && 
b[45650] == 45650 && 
b[45651] == 45651 && 
b[45652] == 45652 && 
b[45653] == 45653 && 
b[45654] == 45654 && 
b[45655] == 45655 && 
b[45656] == 45656 && 
b[45657] == 45657 && 
b[45658] == 45658 && 
b[45659] == 45659 && 
b[45660] == 45660 && 
b[45661] == 45661 && 
b[45662] == 45662 && 
b[45663] == 45663 && 
b[45664] == 45664 && 
b[45665] == 45665 && 
b[45666] == 45666 && 
b[45667] == 45667 && 
b[45668] == 45668 && 
b[45669] == 45669 && 
b[45670] == 45670 && 
b[45671] == 45671 && 
b[45672] == 45672 && 
b[45673] == 45673 && 
b[45674] == 45674 && 
b[45675] == 45675 && 
b[45676] == 45676 && 
b[45677] == 45677 && 
b[45678] == 45678 && 
b[45679] == 45679 && 
b[45680] == 45680 && 
b[45681] == 45681 && 
b[45682] == 45682 && 
b[45683] == 45683 && 
b[45684] == 45684 && 
b[45685] == 45685 && 
b[45686] == 45686 && 
b[45687] == 45687 && 
b[45688] == 45688 && 
b[45689] == 45689 && 
b[45690] == 45690 && 
b[45691] == 45691 && 
b[45692] == 45692 && 
b[45693] == 45693 && 
b[45694] == 45694 && 
b[45695] == 45695 && 
b[45696] == 45696 && 
b[45697] == 45697 && 
b[45698] == 45698 && 
b[45699] == 45699 && 
b[45700] == 45700 && 
b[45701] == 45701 && 
b[45702] == 45702 && 
b[45703] == 45703 && 
b[45704] == 45704 && 
b[45705] == 45705 && 
b[45706] == 45706 && 
b[45707] == 45707 && 
b[45708] == 45708 && 
b[45709] == 45709 && 
b[45710] == 45710 && 
b[45711] == 45711 && 
b[45712] == 45712 && 
b[45713] == 45713 && 
b[45714] == 45714 && 
b[45715] == 45715 && 
b[45716] == 45716 && 
b[45717] == 45717 && 
b[45718] == 45718 && 
b[45719] == 45719 && 
b[45720] == 45720 && 
b[45721] == 45721 && 
b[45722] == 45722 && 
b[45723] == 45723 && 
b[45724] == 45724 && 
b[45725] == 45725 && 
b[45726] == 45726 && 
b[45727] == 45727 && 
b[45728] == 45728 && 
b[45729] == 45729 && 
b[45730] == 45730 && 
b[45731] == 45731 && 
b[45732] == 45732 && 
b[45733] == 45733 && 
b[45734] == 45734 && 
b[45735] == 45735 && 
b[45736] == 45736 && 
b[45737] == 45737 && 
b[45738] == 45738 && 
b[45739] == 45739 && 
b[45740] == 45740 && 
b[45741] == 45741 && 
b[45742] == 45742 && 
b[45743] == 45743 && 
b[45744] == 45744 && 
b[45745] == 45745 && 
b[45746] == 45746 && 
b[45747] == 45747 && 
b[45748] == 45748 && 
b[45749] == 45749 && 
b[45750] == 45750 && 
b[45751] == 45751 && 
b[45752] == 45752 && 
b[45753] == 45753 && 
b[45754] == 45754 && 
b[45755] == 45755 && 
b[45756] == 45756 && 
b[45757] == 45757 && 
b[45758] == 45758 && 
b[45759] == 45759 && 
b[45760] == 45760 && 
b[45761] == 45761 && 
b[45762] == 45762 && 
b[45763] == 45763 && 
b[45764] == 45764 && 
b[45765] == 45765 && 
b[45766] == 45766 && 
b[45767] == 45767 && 
b[45768] == 45768 && 
b[45769] == 45769 && 
b[45770] == 45770 && 
b[45771] == 45771 && 
b[45772] == 45772 && 
b[45773] == 45773 && 
b[45774] == 45774 && 
b[45775] == 45775 && 
b[45776] == 45776 && 
b[45777] == 45777 && 
b[45778] == 45778 && 
b[45779] == 45779 && 
b[45780] == 45780 && 
b[45781] == 45781 && 
b[45782] == 45782 && 
b[45783] == 45783 && 
b[45784] == 45784 && 
b[45785] == 45785 && 
b[45786] == 45786 && 
b[45787] == 45787 && 
b[45788] == 45788 && 
b[45789] == 45789 && 
b[45790] == 45790 && 
b[45791] == 45791 && 
b[45792] == 45792 && 
b[45793] == 45793 && 
b[45794] == 45794 && 
b[45795] == 45795 && 
b[45796] == 45796 && 
b[45797] == 45797 && 
b[45798] == 45798 && 
b[45799] == 45799 && 
b[45800] == 45800 && 
b[45801] == 45801 && 
b[45802] == 45802 && 
b[45803] == 45803 && 
b[45804] == 45804 && 
b[45805] == 45805 && 
b[45806] == 45806 && 
b[45807] == 45807 && 
b[45808] == 45808 && 
b[45809] == 45809 && 
b[45810] == 45810 && 
b[45811] == 45811 && 
b[45812] == 45812 && 
b[45813] == 45813 && 
b[45814] == 45814 && 
b[45815] == 45815 && 
b[45816] == 45816 && 
b[45817] == 45817 && 
b[45818] == 45818 && 
b[45819] == 45819 && 
b[45820] == 45820 && 
b[45821] == 45821 && 
b[45822] == 45822 && 
b[45823] == 45823 && 
b[45824] == 45824 && 
b[45825] == 45825 && 
b[45826] == 45826 && 
b[45827] == 45827 && 
b[45828] == 45828 && 
b[45829] == 45829 && 
b[45830] == 45830 && 
b[45831] == 45831 && 
b[45832] == 45832 && 
b[45833] == 45833 && 
b[45834] == 45834 && 
b[45835] == 45835 && 
b[45836] == 45836 && 
b[45837] == 45837 && 
b[45838] == 45838 && 
b[45839] == 45839 && 
b[45840] == 45840 && 
b[45841] == 45841 && 
b[45842] == 45842 && 
b[45843] == 45843 && 
b[45844] == 45844 && 
b[45845] == 45845 && 
b[45846] == 45846 && 
b[45847] == 45847 && 
b[45848] == 45848 && 
b[45849] == 45849 && 
b[45850] == 45850 && 
b[45851] == 45851 && 
b[45852] == 45852 && 
b[45853] == 45853 && 
b[45854] == 45854 && 
b[45855] == 45855 && 
b[45856] == 45856 && 
b[45857] == 45857 && 
b[45858] == 45858 && 
b[45859] == 45859 && 
b[45860] == 45860 && 
b[45861] == 45861 && 
b[45862] == 45862 && 
b[45863] == 45863 && 
b[45864] == 45864 && 
b[45865] == 45865 && 
b[45866] == 45866 && 
b[45867] == 45867 && 
b[45868] == 45868 && 
b[45869] == 45869 && 
b[45870] == 45870 && 
b[45871] == 45871 && 
b[45872] == 45872 && 
b[45873] == 45873 && 
b[45874] == 45874 && 
b[45875] == 45875 && 
b[45876] == 45876 && 
b[45877] == 45877 && 
b[45878] == 45878 && 
b[45879] == 45879 && 
b[45880] == 45880 && 
b[45881] == 45881 && 
b[45882] == 45882 && 
b[45883] == 45883 && 
b[45884] == 45884 && 
b[45885] == 45885 && 
b[45886] == 45886 && 
b[45887] == 45887 && 
b[45888] == 45888 && 
b[45889] == 45889 && 
b[45890] == 45890 && 
b[45891] == 45891 && 
b[45892] == 45892 && 
b[45893] == 45893 && 
b[45894] == 45894 && 
b[45895] == 45895 && 
b[45896] == 45896 && 
b[45897] == 45897 && 
b[45898] == 45898 && 
b[45899] == 45899 && 
b[45900] == 45900 && 
b[45901] == 45901 && 
b[45902] == 45902 && 
b[45903] == 45903 && 
b[45904] == 45904 && 
b[45905] == 45905 && 
b[45906] == 45906 && 
b[45907] == 45907 && 
b[45908] == 45908 && 
b[45909] == 45909 && 
b[45910] == 45910 && 
b[45911] == 45911 && 
b[45912] == 45912 && 
b[45913] == 45913 && 
b[45914] == 45914 && 
b[45915] == 45915 && 
b[45916] == 45916 && 
b[45917] == 45917 && 
b[45918] == 45918 && 
b[45919] == 45919 && 
b[45920] == 45920 && 
b[45921] == 45921 && 
b[45922] == 45922 && 
b[45923] == 45923 && 
b[45924] == 45924 && 
b[45925] == 45925 && 
b[45926] == 45926 && 
b[45927] == 45927 && 
b[45928] == 45928 && 
b[45929] == 45929 && 
b[45930] == 45930 && 
b[45931] == 45931 && 
b[45932] == 45932 && 
b[45933] == 45933 && 
b[45934] == 45934 && 
b[45935] == 45935 && 
b[45936] == 45936 && 
b[45937] == 45937 && 
b[45938] == 45938 && 
b[45939] == 45939 && 
b[45940] == 45940 && 
b[45941] == 45941 && 
b[45942] == 45942 && 
b[45943] == 45943 && 
b[45944] == 45944 && 
b[45945] == 45945 && 
b[45946] == 45946 && 
b[45947] == 45947 && 
b[45948] == 45948 && 
b[45949] == 45949 && 
b[45950] == 45950 && 
b[45951] == 45951 && 
b[45952] == 45952 && 
b[45953] == 45953 && 
b[45954] == 45954 && 
b[45955] == 45955 && 
b[45956] == 45956 && 
b[45957] == 45957 && 
b[45958] == 45958 && 
b[45959] == 45959 && 
b[45960] == 45960 && 
b[45961] == 45961 && 
b[45962] == 45962 && 
b[45963] == 45963 && 
b[45964] == 45964 && 
b[45965] == 45965 && 
b[45966] == 45966 && 
b[45967] == 45967 && 
b[45968] == 45968 && 
b[45969] == 45969 && 
b[45970] == 45970 && 
b[45971] == 45971 && 
b[45972] == 45972 && 
b[45973] == 45973 && 
b[45974] == 45974 && 
b[45975] == 45975 && 
b[45976] == 45976 && 
b[45977] == 45977 && 
b[45978] == 45978 && 
b[45979] == 45979 && 
b[45980] == 45980 && 
b[45981] == 45981 && 
b[45982] == 45982 && 
b[45983] == 45983 && 
b[45984] == 45984 && 
b[45985] == 45985 && 
b[45986] == 45986 && 
b[45987] == 45987 && 
b[45988] == 45988 && 
b[45989] == 45989 && 
b[45990] == 45990 && 
b[45991] == 45991 && 
b[45992] == 45992 && 
b[45993] == 45993 && 
b[45994] == 45994 && 
b[45995] == 45995 && 
b[45996] == 45996 && 
b[45997] == 45997 && 
b[45998] == 45998 && 
b[45999] == 45999 && 
b[46000] == 46000 && 
b[46001] == 46001 && 
b[46002] == 46002 && 
b[46003] == 46003 && 
b[46004] == 46004 && 
b[46005] == 46005 && 
b[46006] == 46006 && 
b[46007] == 46007 && 
b[46008] == 46008 && 
b[46009] == 46009 && 
b[46010] == 46010 && 
b[46011] == 46011 && 
b[46012] == 46012 && 
b[46013] == 46013 && 
b[46014] == 46014 && 
b[46015] == 46015 && 
b[46016] == 46016 && 
b[46017] == 46017 && 
b[46018] == 46018 && 
b[46019] == 46019 && 
b[46020] == 46020 && 
b[46021] == 46021 && 
b[46022] == 46022 && 
b[46023] == 46023 && 
b[46024] == 46024 && 
b[46025] == 46025 && 
b[46026] == 46026 && 
b[46027] == 46027 && 
b[46028] == 46028 && 
b[46029] == 46029 && 
b[46030] == 46030 && 
b[46031] == 46031 && 
b[46032] == 46032 && 
b[46033] == 46033 && 
b[46034] == 46034 && 
b[46035] == 46035 && 
b[46036] == 46036 && 
b[46037] == 46037 && 
b[46038] == 46038 && 
b[46039] == 46039 && 
b[46040] == 46040 && 
b[46041] == 46041 && 
b[46042] == 46042 && 
b[46043] == 46043 && 
b[46044] == 46044 && 
b[46045] == 46045 && 
b[46046] == 46046 && 
b[46047] == 46047 && 
b[46048] == 46048 && 
b[46049] == 46049 && 
b[46050] == 46050 && 
b[46051] == 46051 && 
b[46052] == 46052 && 
b[46053] == 46053 && 
b[46054] == 46054 && 
b[46055] == 46055 && 
b[46056] == 46056 && 
b[46057] == 46057 && 
b[46058] == 46058 && 
b[46059] == 46059 && 
b[46060] == 46060 && 
b[46061] == 46061 && 
b[46062] == 46062 && 
b[46063] == 46063 && 
b[46064] == 46064 && 
b[46065] == 46065 && 
b[46066] == 46066 && 
b[46067] == 46067 && 
b[46068] == 46068 && 
b[46069] == 46069 && 
b[46070] == 46070 && 
b[46071] == 46071 && 
b[46072] == 46072 && 
b[46073] == 46073 && 
b[46074] == 46074 && 
b[46075] == 46075 && 
b[46076] == 46076 && 
b[46077] == 46077 && 
b[46078] == 46078 && 
b[46079] == 46079 && 
b[46080] == 46080 && 
b[46081] == 46081 && 
b[46082] == 46082 && 
b[46083] == 46083 && 
b[46084] == 46084 && 
b[46085] == 46085 && 
b[46086] == 46086 && 
b[46087] == 46087 && 
b[46088] == 46088 && 
b[46089] == 46089 && 
b[46090] == 46090 && 
b[46091] == 46091 && 
b[46092] == 46092 && 
b[46093] == 46093 && 
b[46094] == 46094 && 
b[46095] == 46095 && 
b[46096] == 46096 && 
b[46097] == 46097 && 
b[46098] == 46098 && 
b[46099] == 46099 && 
b[46100] == 46100 && 
b[46101] == 46101 && 
b[46102] == 46102 && 
b[46103] == 46103 && 
b[46104] == 46104 && 
b[46105] == 46105 && 
b[46106] == 46106 && 
b[46107] == 46107 && 
b[46108] == 46108 && 
b[46109] == 46109 && 
b[46110] == 46110 && 
b[46111] == 46111 && 
b[46112] == 46112 && 
b[46113] == 46113 && 
b[46114] == 46114 && 
b[46115] == 46115 && 
b[46116] == 46116 && 
b[46117] == 46117 && 
b[46118] == 46118 && 
b[46119] == 46119 && 
b[46120] == 46120 && 
b[46121] == 46121 && 
b[46122] == 46122 && 
b[46123] == 46123 && 
b[46124] == 46124 && 
b[46125] == 46125 && 
b[46126] == 46126 && 
b[46127] == 46127 && 
b[46128] == 46128 && 
b[46129] == 46129 && 
b[46130] == 46130 && 
b[46131] == 46131 && 
b[46132] == 46132 && 
b[46133] == 46133 && 
b[46134] == 46134 && 
b[46135] == 46135 && 
b[46136] == 46136 && 
b[46137] == 46137 && 
b[46138] == 46138 && 
b[46139] == 46139 && 
b[46140] == 46140 && 
b[46141] == 46141 && 
b[46142] == 46142 && 
b[46143] == 46143 && 
b[46144] == 46144 && 
b[46145] == 46145 && 
b[46146] == 46146 && 
b[46147] == 46147 && 
b[46148] == 46148 && 
b[46149] == 46149 && 
b[46150] == 46150 && 
b[46151] == 46151 && 
b[46152] == 46152 && 
b[46153] == 46153 && 
b[46154] == 46154 && 
b[46155] == 46155 && 
b[46156] == 46156 && 
b[46157] == 46157 && 
b[46158] == 46158 && 
b[46159] == 46159 && 
b[46160] == 46160 && 
b[46161] == 46161 && 
b[46162] == 46162 && 
b[46163] == 46163 && 
b[46164] == 46164 && 
b[46165] == 46165 && 
b[46166] == 46166 && 
b[46167] == 46167 && 
b[46168] == 46168 && 
b[46169] == 46169 && 
b[46170] == 46170 && 
b[46171] == 46171 && 
b[46172] == 46172 && 
b[46173] == 46173 && 
b[46174] == 46174 && 
b[46175] == 46175 && 
b[46176] == 46176 && 
b[46177] == 46177 && 
b[46178] == 46178 && 
b[46179] == 46179 && 
b[46180] == 46180 && 
b[46181] == 46181 && 
b[46182] == 46182 && 
b[46183] == 46183 && 
b[46184] == 46184 && 
b[46185] == 46185 && 
b[46186] == 46186 && 
b[46187] == 46187 && 
b[46188] == 46188 && 
b[46189] == 46189 && 
b[46190] == 46190 && 
b[46191] == 46191 && 
b[46192] == 46192 && 
b[46193] == 46193 && 
b[46194] == 46194 && 
b[46195] == 46195 && 
b[46196] == 46196 && 
b[46197] == 46197 && 
b[46198] == 46198 && 
b[46199] == 46199 && 
b[46200] == 46200 && 
b[46201] == 46201 && 
b[46202] == 46202 && 
b[46203] == 46203 && 
b[46204] == 46204 && 
b[46205] == 46205 && 
b[46206] == 46206 && 
b[46207] == 46207 && 
b[46208] == 46208 && 
b[46209] == 46209 && 
b[46210] == 46210 && 
b[46211] == 46211 && 
b[46212] == 46212 && 
b[46213] == 46213 && 
b[46214] == 46214 && 
b[46215] == 46215 && 
b[46216] == 46216 && 
b[46217] == 46217 && 
b[46218] == 46218 && 
b[46219] == 46219 && 
b[46220] == 46220 && 
b[46221] == 46221 && 
b[46222] == 46222 && 
b[46223] == 46223 && 
b[46224] == 46224 && 
b[46225] == 46225 && 
b[46226] == 46226 && 
b[46227] == 46227 && 
b[46228] == 46228 && 
b[46229] == 46229 && 
b[46230] == 46230 && 
b[46231] == 46231 && 
b[46232] == 46232 && 
b[46233] == 46233 && 
b[46234] == 46234 && 
b[46235] == 46235 && 
b[46236] == 46236 && 
b[46237] == 46237 && 
b[46238] == 46238 && 
b[46239] == 46239 && 
b[46240] == 46240 && 
b[46241] == 46241 && 
b[46242] == 46242 && 
b[46243] == 46243 && 
b[46244] == 46244 && 
b[46245] == 46245 && 
b[46246] == 46246 && 
b[46247] == 46247 && 
b[46248] == 46248 && 
b[46249] == 46249 && 
b[46250] == 46250 && 
b[46251] == 46251 && 
b[46252] == 46252 && 
b[46253] == 46253 && 
b[46254] == 46254 && 
b[46255] == 46255 && 
b[46256] == 46256 && 
b[46257] == 46257 && 
b[46258] == 46258 && 
b[46259] == 46259 && 
b[46260] == 46260 && 
b[46261] == 46261 && 
b[46262] == 46262 && 
b[46263] == 46263 && 
b[46264] == 46264 && 
b[46265] == 46265 && 
b[46266] == 46266 && 
b[46267] == 46267 && 
b[46268] == 46268 && 
b[46269] == 46269 && 
b[46270] == 46270 && 
b[46271] == 46271 && 
b[46272] == 46272 && 
b[46273] == 46273 && 
b[46274] == 46274 && 
b[46275] == 46275 && 
b[46276] == 46276 && 
b[46277] == 46277 && 
b[46278] == 46278 && 
b[46279] == 46279 && 
b[46280] == 46280 && 
b[46281] == 46281 && 
b[46282] == 46282 && 
b[46283] == 46283 && 
b[46284] == 46284 && 
b[46285] == 46285 && 
b[46286] == 46286 && 
b[46287] == 46287 && 
b[46288] == 46288 && 
b[46289] == 46289 && 
b[46290] == 46290 && 
b[46291] == 46291 && 
b[46292] == 46292 && 
b[46293] == 46293 && 
b[46294] == 46294 && 
b[46295] == 46295 && 
b[46296] == 46296 && 
b[46297] == 46297 && 
b[46298] == 46298 && 
b[46299] == 46299 && 
b[46300] == 46300 && 
b[46301] == 46301 && 
b[46302] == 46302 && 
b[46303] == 46303 && 
b[46304] == 46304 && 
b[46305] == 46305 && 
b[46306] == 46306 && 
b[46307] == 46307 && 
b[46308] == 46308 && 
b[46309] == 46309 && 
b[46310] == 46310 && 
b[46311] == 46311 && 
b[46312] == 46312 && 
b[46313] == 46313 && 
b[46314] == 46314 && 
b[46315] == 46315 && 
b[46316] == 46316 && 
b[46317] == 46317 && 
b[46318] == 46318 && 
b[46319] == 46319 && 
b[46320] == 46320 && 
b[46321] == 46321 && 
b[46322] == 46322 && 
b[46323] == 46323 && 
b[46324] == 46324 && 
b[46325] == 46325 && 
b[46326] == 46326 && 
b[46327] == 46327 && 
b[46328] == 46328 && 
b[46329] == 46329 && 
b[46330] == 46330 && 
b[46331] == 46331 && 
b[46332] == 46332 && 
b[46333] == 46333 && 
b[46334] == 46334 && 
b[46335] == 46335 && 
b[46336] == 46336 && 
b[46337] == 46337 && 
b[46338] == 46338 && 
b[46339] == 46339 && 
b[46340] == 46340 && 
b[46341] == 46341 && 
b[46342] == 46342 && 
b[46343] == 46343 && 
b[46344] == 46344 && 
b[46345] == 46345 && 
b[46346] == 46346 && 
b[46347] == 46347 && 
b[46348] == 46348 && 
b[46349] == 46349 && 
b[46350] == 46350 && 
b[46351] == 46351 && 
b[46352] == 46352 && 
b[46353] == 46353 && 
b[46354] == 46354 && 
b[46355] == 46355 && 
b[46356] == 46356 && 
b[46357] == 46357 && 
b[46358] == 46358 && 
b[46359] == 46359 && 
b[46360] == 46360 && 
b[46361] == 46361 && 
b[46362] == 46362 && 
b[46363] == 46363 && 
b[46364] == 46364 && 
b[46365] == 46365 && 
b[46366] == 46366 && 
b[46367] == 46367 && 
b[46368] == 46368 && 
b[46369] == 46369 && 
b[46370] == 46370 && 
b[46371] == 46371 && 
b[46372] == 46372 && 
b[46373] == 46373 && 
b[46374] == 46374 && 
b[46375] == 46375 && 
b[46376] == 46376 && 
b[46377] == 46377 && 
b[46378] == 46378 && 
b[46379] == 46379 && 
b[46380] == 46380 && 
b[46381] == 46381 && 
b[46382] == 46382 && 
b[46383] == 46383 && 
b[46384] == 46384 && 
b[46385] == 46385 && 
b[46386] == 46386 && 
b[46387] == 46387 && 
b[46388] == 46388 && 
b[46389] == 46389 && 
b[46390] == 46390 && 
b[46391] == 46391 && 
b[46392] == 46392 && 
b[46393] == 46393 && 
b[46394] == 46394 && 
b[46395] == 46395 && 
b[46396] == 46396 && 
b[46397] == 46397 && 
b[46398] == 46398 && 
b[46399] == 46399 && 
b[46400] == 46400 && 
b[46401] == 46401 && 
b[46402] == 46402 && 
b[46403] == 46403 && 
b[46404] == 46404 && 
b[46405] == 46405 && 
b[46406] == 46406 && 
b[46407] == 46407 && 
b[46408] == 46408 && 
b[46409] == 46409 && 
b[46410] == 46410 && 
b[46411] == 46411 && 
b[46412] == 46412 && 
b[46413] == 46413 && 
b[46414] == 46414 && 
b[46415] == 46415 && 
b[46416] == 46416 && 
b[46417] == 46417 && 
b[46418] == 46418 && 
b[46419] == 46419 && 
b[46420] == 46420 && 
b[46421] == 46421 && 
b[46422] == 46422 && 
b[46423] == 46423 && 
b[46424] == 46424 && 
b[46425] == 46425 && 
b[46426] == 46426 && 
b[46427] == 46427 && 
b[46428] == 46428 && 
b[46429] == 46429 && 
b[46430] == 46430 && 
b[46431] == 46431 && 
b[46432] == 46432 && 
b[46433] == 46433 && 
b[46434] == 46434 && 
b[46435] == 46435 && 
b[46436] == 46436 && 
b[46437] == 46437 && 
b[46438] == 46438 && 
b[46439] == 46439 && 
b[46440] == 46440 && 
b[46441] == 46441 && 
b[46442] == 46442 && 
b[46443] == 46443 && 
b[46444] == 46444 && 
b[46445] == 46445 && 
b[46446] == 46446 && 
b[46447] == 46447 && 
b[46448] == 46448 && 
b[46449] == 46449 && 
b[46450] == 46450 && 
b[46451] == 46451 && 
b[46452] == 46452 && 
b[46453] == 46453 && 
b[46454] == 46454 && 
b[46455] == 46455 && 
b[46456] == 46456 && 
b[46457] == 46457 && 
b[46458] == 46458 && 
b[46459] == 46459 && 
b[46460] == 46460 && 
b[46461] == 46461 && 
b[46462] == 46462 && 
b[46463] == 46463 && 
b[46464] == 46464 && 
b[46465] == 46465 && 
b[46466] == 46466 && 
b[46467] == 46467 && 
b[46468] == 46468 && 
b[46469] == 46469 && 
b[46470] == 46470 && 
b[46471] == 46471 && 
b[46472] == 46472 && 
b[46473] == 46473 && 
b[46474] == 46474 && 
b[46475] == 46475 && 
b[46476] == 46476 && 
b[46477] == 46477 && 
b[46478] == 46478 && 
b[46479] == 46479 && 
b[46480] == 46480 && 
b[46481] == 46481 && 
b[46482] == 46482 && 
b[46483] == 46483 && 
b[46484] == 46484 && 
b[46485] == 46485 && 
b[46486] == 46486 && 
b[46487] == 46487 && 
b[46488] == 46488 && 
b[46489] == 46489 && 
b[46490] == 46490 && 
b[46491] == 46491 && 
b[46492] == 46492 && 
b[46493] == 46493 && 
b[46494] == 46494 && 
b[46495] == 46495 && 
b[46496] == 46496 && 
b[46497] == 46497 && 
b[46498] == 46498 && 
b[46499] == 46499 && 
b[46500] == 46500 && 
b[46501] == 46501 && 
b[46502] == 46502 && 
b[46503] == 46503 && 
b[46504] == 46504 && 
b[46505] == 46505 && 
b[46506] == 46506 && 
b[46507] == 46507 && 
b[46508] == 46508 && 
b[46509] == 46509 && 
b[46510] == 46510 && 
b[46511] == 46511 && 
b[46512] == 46512 && 
b[46513] == 46513 && 
b[46514] == 46514 && 
b[46515] == 46515 && 
b[46516] == 46516 && 
b[46517] == 46517 && 
b[46518] == 46518 && 
b[46519] == 46519 && 
b[46520] == 46520 && 
b[46521] == 46521 && 
b[46522] == 46522 && 
b[46523] == 46523 && 
b[46524] == 46524 && 
b[46525] == 46525 && 
b[46526] == 46526 && 
b[46527] == 46527 && 
b[46528] == 46528 && 
b[46529] == 46529 && 
b[46530] == 46530 && 
b[46531] == 46531 && 
b[46532] == 46532 && 
b[46533] == 46533 && 
b[46534] == 46534 && 
b[46535] == 46535 && 
b[46536] == 46536 && 
b[46537] == 46537 && 
b[46538] == 46538 && 
b[46539] == 46539 && 
b[46540] == 46540 && 
b[46541] == 46541 && 
b[46542] == 46542 && 
b[46543] == 46543 && 
b[46544] == 46544 && 
b[46545] == 46545 && 
b[46546] == 46546 && 
b[46547] == 46547 && 
b[46548] == 46548 && 
b[46549] == 46549 && 
b[46550] == 46550 && 
b[46551] == 46551 && 
b[46552] == 46552 && 
b[46553] == 46553 && 
b[46554] == 46554 && 
b[46555] == 46555 && 
b[46556] == 46556 && 
b[46557] == 46557 && 
b[46558] == 46558 && 
b[46559] == 46559 && 
b[46560] == 46560 && 
b[46561] == 46561 && 
b[46562] == 46562 && 
b[46563] == 46563 && 
b[46564] == 46564 && 
b[46565] == 46565 && 
b[46566] == 46566 && 
b[46567] == 46567 && 
b[46568] == 46568 && 
b[46569] == 46569 && 
b[46570] == 46570 && 
b[46571] == 46571 && 
b[46572] == 46572 && 
b[46573] == 46573 && 
b[46574] == 46574 && 
b[46575] == 46575 && 
b[46576] == 46576 && 
b[46577] == 46577 && 
b[46578] == 46578 && 
b[46579] == 46579 && 
b[46580] == 46580 && 
b[46581] == 46581 && 
b[46582] == 46582 && 
b[46583] == 46583 && 
b[46584] == 46584 && 
b[46585] == 46585 && 
b[46586] == 46586 && 
b[46587] == 46587 && 
b[46588] == 46588 && 
b[46589] == 46589 && 
b[46590] == 46590 && 
b[46591] == 46591 && 
b[46592] == 46592 && 
b[46593] == 46593 && 
b[46594] == 46594 && 
b[46595] == 46595 && 
b[46596] == 46596 && 
b[46597] == 46597 && 
b[46598] == 46598 && 
b[46599] == 46599 && 
b[46600] == 46600 && 
b[46601] == 46601 && 
b[46602] == 46602 && 
b[46603] == 46603 && 
b[46604] == 46604 && 
b[46605] == 46605 && 
b[46606] == 46606 && 
b[46607] == 46607 && 
b[46608] == 46608 && 
b[46609] == 46609 && 
b[46610] == 46610 && 
b[46611] == 46611 && 
b[46612] == 46612 && 
b[46613] == 46613 && 
b[46614] == 46614 && 
b[46615] == 46615 && 
b[46616] == 46616 && 
b[46617] == 46617 && 
b[46618] == 46618 && 
b[46619] == 46619 && 
b[46620] == 46620 && 
b[46621] == 46621 && 
b[46622] == 46622 && 
b[46623] == 46623 && 
b[46624] == 46624 && 
b[46625] == 46625 && 
b[46626] == 46626 && 
b[46627] == 46627 && 
b[46628] == 46628 && 
b[46629] == 46629 && 
b[46630] == 46630 && 
b[46631] == 46631 && 
b[46632] == 46632 && 
b[46633] == 46633 && 
b[46634] == 46634 && 
b[46635] == 46635 && 
b[46636] == 46636 && 
b[46637] == 46637 && 
b[46638] == 46638 && 
b[46639] == 46639 && 
b[46640] == 46640 && 
b[46641] == 46641 && 
b[46642] == 46642 && 
b[46643] == 46643 && 
b[46644] == 46644 && 
b[46645] == 46645 && 
b[46646] == 46646 && 
b[46647] == 46647 && 
b[46648] == 46648 && 
b[46649] == 46649 && 
b[46650] == 46650 && 
b[46651] == 46651 && 
b[46652] == 46652 && 
b[46653] == 46653 && 
b[46654] == 46654 && 
b[46655] == 46655 && 
b[46656] == 46656 && 
b[46657] == 46657 && 
b[46658] == 46658 && 
b[46659] == 46659 && 
b[46660] == 46660 && 
b[46661] == 46661 && 
b[46662] == 46662 && 
b[46663] == 46663 && 
b[46664] == 46664 && 
b[46665] == 46665 && 
b[46666] == 46666 && 
b[46667] == 46667 && 
b[46668] == 46668 && 
b[46669] == 46669 && 
b[46670] == 46670 && 
b[46671] == 46671 && 
b[46672] == 46672 && 
b[46673] == 46673 && 
b[46674] == 46674 && 
b[46675] == 46675 && 
b[46676] == 46676 && 
b[46677] == 46677 && 
b[46678] == 46678 && 
b[46679] == 46679 && 
b[46680] == 46680 && 
b[46681] == 46681 && 
b[46682] == 46682 && 
b[46683] == 46683 && 
b[46684] == 46684 && 
b[46685] == 46685 && 
b[46686] == 46686 && 
b[46687] == 46687 && 
b[46688] == 46688 && 
b[46689] == 46689 && 
b[46690] == 46690 && 
b[46691] == 46691 && 
b[46692] == 46692 && 
b[46693] == 46693 && 
b[46694] == 46694 && 
b[46695] == 46695 && 
b[46696] == 46696 && 
b[46697] == 46697 && 
b[46698] == 46698 && 
b[46699] == 46699 && 
b[46700] == 46700 && 
b[46701] == 46701 && 
b[46702] == 46702 && 
b[46703] == 46703 && 
b[46704] == 46704 && 
b[46705] == 46705 && 
b[46706] == 46706 && 
b[46707] == 46707 && 
b[46708] == 46708 && 
b[46709] == 46709 && 
b[46710] == 46710 && 
b[46711] == 46711 && 
b[46712] == 46712 && 
b[46713] == 46713 && 
b[46714] == 46714 && 
b[46715] == 46715 && 
b[46716] == 46716 && 
b[46717] == 46717 && 
b[46718] == 46718 && 
b[46719] == 46719 && 
b[46720] == 46720 && 
b[46721] == 46721 && 
b[46722] == 46722 && 
b[46723] == 46723 && 
b[46724] == 46724 && 
b[46725] == 46725 && 
b[46726] == 46726 && 
b[46727] == 46727 && 
b[46728] == 46728 && 
b[46729] == 46729 && 
b[46730] == 46730 && 
b[46731] == 46731 && 
b[46732] == 46732 && 
b[46733] == 46733 && 
b[46734] == 46734 && 
b[46735] == 46735 && 
b[46736] == 46736 && 
b[46737] == 46737 && 
b[46738] == 46738 && 
b[46739] == 46739 && 
b[46740] == 46740 && 
b[46741] == 46741 && 
b[46742] == 46742 && 
b[46743] == 46743 && 
b[46744] == 46744 && 
b[46745] == 46745 && 
b[46746] == 46746 && 
b[46747] == 46747 && 
b[46748] == 46748 && 
b[46749] == 46749 && 
b[46750] == 46750 && 
b[46751] == 46751 && 
b[46752] == 46752 && 
b[46753] == 46753 && 
b[46754] == 46754 && 
b[46755] == 46755 && 
b[46756] == 46756 && 
b[46757] == 46757 && 
b[46758] == 46758 && 
b[46759] == 46759 && 
b[46760] == 46760 && 
b[46761] == 46761 && 
b[46762] == 46762 && 
b[46763] == 46763 && 
b[46764] == 46764 && 
b[46765] == 46765 && 
b[46766] == 46766 && 
b[46767] == 46767 && 
b[46768] == 46768 && 
b[46769] == 46769 && 
b[46770] == 46770 && 
b[46771] == 46771 && 
b[46772] == 46772 && 
b[46773] == 46773 && 
b[46774] == 46774 && 
b[46775] == 46775 && 
b[46776] == 46776 && 
b[46777] == 46777 && 
b[46778] == 46778 && 
b[46779] == 46779 && 
b[46780] == 46780 && 
b[46781] == 46781 && 
b[46782] == 46782 && 
b[46783] == 46783 && 
b[46784] == 46784 && 
b[46785] == 46785 && 
b[46786] == 46786 && 
b[46787] == 46787 && 
b[46788] == 46788 && 
b[46789] == 46789 && 
b[46790] == 46790 && 
b[46791] == 46791 && 
b[46792] == 46792 && 
b[46793] == 46793 && 
b[46794] == 46794 && 
b[46795] == 46795 && 
b[46796] == 46796 && 
b[46797] == 46797 && 
b[46798] == 46798 && 
b[46799] == 46799 && 
b[46800] == 46800 && 
b[46801] == 46801 && 
b[46802] == 46802 && 
b[46803] == 46803 && 
b[46804] == 46804 && 
b[46805] == 46805 && 
b[46806] == 46806 && 
b[46807] == 46807 && 
b[46808] == 46808 && 
b[46809] == 46809 && 
b[46810] == 46810 && 
b[46811] == 46811 && 
b[46812] == 46812 && 
b[46813] == 46813 && 
b[46814] == 46814 && 
b[46815] == 46815 && 
b[46816] == 46816 && 
b[46817] == 46817 && 
b[46818] == 46818 && 
b[46819] == 46819 && 
b[46820] == 46820 && 
b[46821] == 46821 && 
b[46822] == 46822 && 
b[46823] == 46823 && 
b[46824] == 46824 && 
b[46825] == 46825 && 
b[46826] == 46826 && 
b[46827] == 46827 && 
b[46828] == 46828 && 
b[46829] == 46829 && 
b[46830] == 46830 && 
b[46831] == 46831 && 
b[46832] == 46832 && 
b[46833] == 46833 && 
b[46834] == 46834 && 
b[46835] == 46835 && 
b[46836] == 46836 && 
b[46837] == 46837 && 
b[46838] == 46838 && 
b[46839] == 46839 && 
b[46840] == 46840 && 
b[46841] == 46841 && 
b[46842] == 46842 && 
b[46843] == 46843 && 
b[46844] == 46844 && 
b[46845] == 46845 && 
b[46846] == 46846 && 
b[46847] == 46847 && 
b[46848] == 46848 && 
b[46849] == 46849 && 
b[46850] == 46850 && 
b[46851] == 46851 && 
b[46852] == 46852 && 
b[46853] == 46853 && 
b[46854] == 46854 && 
b[46855] == 46855 && 
b[46856] == 46856 && 
b[46857] == 46857 && 
b[46858] == 46858 && 
b[46859] == 46859 && 
b[46860] == 46860 && 
b[46861] == 46861 && 
b[46862] == 46862 && 
b[46863] == 46863 && 
b[46864] == 46864 && 
b[46865] == 46865 && 
b[46866] == 46866 && 
b[46867] == 46867 && 
b[46868] == 46868 && 
b[46869] == 46869 && 
b[46870] == 46870 && 
b[46871] == 46871 && 
b[46872] == 46872 && 
b[46873] == 46873 && 
b[46874] == 46874 && 
b[46875] == 46875 && 
b[46876] == 46876 && 
b[46877] == 46877 && 
b[46878] == 46878 && 
b[46879] == 46879 && 
b[46880] == 46880 && 
b[46881] == 46881 && 
b[46882] == 46882 && 
b[46883] == 46883 && 
b[46884] == 46884 && 
b[46885] == 46885 && 
b[46886] == 46886 && 
b[46887] == 46887 && 
b[46888] == 46888 && 
b[46889] == 46889 && 
b[46890] == 46890 && 
b[46891] == 46891 && 
b[46892] == 46892 && 
b[46893] == 46893 && 
b[46894] == 46894 && 
b[46895] == 46895 && 
b[46896] == 46896 && 
b[46897] == 46897 && 
b[46898] == 46898 && 
b[46899] == 46899 && 
b[46900] == 46900 && 
b[46901] == 46901 && 
b[46902] == 46902 && 
b[46903] == 46903 && 
b[46904] == 46904 && 
b[46905] == 46905 && 
b[46906] == 46906 && 
b[46907] == 46907 && 
b[46908] == 46908 && 
b[46909] == 46909 && 
b[46910] == 46910 && 
b[46911] == 46911 && 
b[46912] == 46912 && 
b[46913] == 46913 && 
b[46914] == 46914 && 
b[46915] == 46915 && 
b[46916] == 46916 && 
b[46917] == 46917 && 
b[46918] == 46918 && 
b[46919] == 46919 && 
b[46920] == 46920 && 
b[46921] == 46921 && 
b[46922] == 46922 && 
b[46923] == 46923 && 
b[46924] == 46924 && 
b[46925] == 46925 && 
b[46926] == 46926 && 
b[46927] == 46927 && 
b[46928] == 46928 && 
b[46929] == 46929 && 
b[46930] == 46930 && 
b[46931] == 46931 && 
b[46932] == 46932 && 
b[46933] == 46933 && 
b[46934] == 46934 && 
b[46935] == 46935 && 
b[46936] == 46936 && 
b[46937] == 46937 && 
b[46938] == 46938 && 
b[46939] == 46939 && 
b[46940] == 46940 && 
b[46941] == 46941 && 
b[46942] == 46942 && 
b[46943] == 46943 && 
b[46944] == 46944 && 
b[46945] == 46945 && 
b[46946] == 46946 && 
b[46947] == 46947 && 
b[46948] == 46948 && 
b[46949] == 46949 && 
b[46950] == 46950 && 
b[46951] == 46951 && 
b[46952] == 46952 && 
b[46953] == 46953 && 
b[46954] == 46954 && 
b[46955] == 46955 && 
b[46956] == 46956 && 
b[46957] == 46957 && 
b[46958] == 46958 && 
b[46959] == 46959 && 
b[46960] == 46960 && 
b[46961] == 46961 && 
b[46962] == 46962 && 
b[46963] == 46963 && 
b[46964] == 46964 && 
b[46965] == 46965 && 
b[46966] == 46966 && 
b[46967] == 46967 && 
b[46968] == 46968 && 
b[46969] == 46969 && 
b[46970] == 46970 && 
b[46971] == 46971 && 
b[46972] == 46972 && 
b[46973] == 46973 && 
b[46974] == 46974 && 
b[46975] == 46975 && 
b[46976] == 46976 && 
b[46977] == 46977 && 
b[46978] == 46978 && 
b[46979] == 46979 && 
b[46980] == 46980 && 
b[46981] == 46981 && 
b[46982] == 46982 && 
b[46983] == 46983 && 
b[46984] == 46984 && 
b[46985] == 46985 && 
b[46986] == 46986 && 
b[46987] == 46987 && 
b[46988] == 46988 && 
b[46989] == 46989 && 
b[46990] == 46990 && 
b[46991] == 46991 && 
b[46992] == 46992 && 
b[46993] == 46993 && 
b[46994] == 46994 && 
b[46995] == 46995 && 
b[46996] == 46996 && 
b[46997] == 46997 && 
b[46998] == 46998 && 
b[46999] == 46999 && 
b[47000] == 47000 && 
b[47001] == 47001 && 
b[47002] == 47002 && 
b[47003] == 47003 && 
b[47004] == 47004 && 
b[47005] == 47005 && 
b[47006] == 47006 && 
b[47007] == 47007 && 
b[47008] == 47008 && 
b[47009] == 47009 && 
b[47010] == 47010 && 
b[47011] == 47011 && 
b[47012] == 47012 && 
b[47013] == 47013 && 
b[47014] == 47014 && 
b[47015] == 47015 && 
b[47016] == 47016 && 
b[47017] == 47017 && 
b[47018] == 47018 && 
b[47019] == 47019 && 
b[47020] == 47020 && 
b[47021] == 47021 && 
b[47022] == 47022 && 
b[47023] == 47023 && 
b[47024] == 47024 && 
b[47025] == 47025 && 
b[47026] == 47026 && 
b[47027] == 47027 && 
b[47028] == 47028 && 
b[47029] == 47029 && 
b[47030] == 47030 && 
b[47031] == 47031 && 
b[47032] == 47032 && 
b[47033] == 47033 && 
b[47034] == 47034 && 
b[47035] == 47035 && 
b[47036] == 47036 && 
b[47037] == 47037 && 
b[47038] == 47038 && 
b[47039] == 47039 && 
b[47040] == 47040 && 
b[47041] == 47041 && 
b[47042] == 47042 && 
b[47043] == 47043 && 
b[47044] == 47044 && 
b[47045] == 47045 && 
b[47046] == 47046 && 
b[47047] == 47047 && 
b[47048] == 47048 && 
b[47049] == 47049 && 
b[47050] == 47050 && 
b[47051] == 47051 && 
b[47052] == 47052 && 
b[47053] == 47053 && 
b[47054] == 47054 && 
b[47055] == 47055 && 
b[47056] == 47056 && 
b[47057] == 47057 && 
b[47058] == 47058 && 
b[47059] == 47059 && 
b[47060] == 47060 && 
b[47061] == 47061 && 
b[47062] == 47062 && 
b[47063] == 47063 && 
b[47064] == 47064 && 
b[47065] == 47065 && 
b[47066] == 47066 && 
b[47067] == 47067 && 
b[47068] == 47068 && 
b[47069] == 47069 && 
b[47070] == 47070 && 
b[47071] == 47071 && 
b[47072] == 47072 && 
b[47073] == 47073 && 
b[47074] == 47074 && 
b[47075] == 47075 && 
b[47076] == 47076 && 
b[47077] == 47077 && 
b[47078] == 47078 && 
b[47079] == 47079 && 
b[47080] == 47080 && 
b[47081] == 47081 && 
b[47082] == 47082 && 
b[47083] == 47083 && 
b[47084] == 47084 && 
b[47085] == 47085 && 
b[47086] == 47086 && 
b[47087] == 47087 && 
b[47088] == 47088 && 
b[47089] == 47089 && 
b[47090] == 47090 && 
b[47091] == 47091 && 
b[47092] == 47092 && 
b[47093] == 47093 && 
b[47094] == 47094 && 
b[47095] == 47095 && 
b[47096] == 47096 && 
b[47097] == 47097 && 
b[47098] == 47098 && 
b[47099] == 47099 && 
b[47100] == 47100 && 
b[47101] == 47101 && 
b[47102] == 47102 && 
b[47103] == 47103 && 
b[47104] == 47104 && 
b[47105] == 47105 && 
b[47106] == 47106 && 
b[47107] == 47107 && 
b[47108] == 47108 && 
b[47109] == 47109 && 
b[47110] == 47110 && 
b[47111] == 47111 && 
b[47112] == 47112 && 
b[47113] == 47113 && 
b[47114] == 47114 && 
b[47115] == 47115 && 
b[47116] == 47116 && 
b[47117] == 47117 && 
b[47118] == 47118 && 
b[47119] == 47119 && 
b[47120] == 47120 && 
b[47121] == 47121 && 
b[47122] == 47122 && 
b[47123] == 47123 && 
b[47124] == 47124 && 
b[47125] == 47125 && 
b[47126] == 47126 && 
b[47127] == 47127 && 
b[47128] == 47128 && 
b[47129] == 47129 && 
b[47130] == 47130 && 
b[47131] == 47131 && 
b[47132] == 47132 && 
b[47133] == 47133 && 
b[47134] == 47134 && 
b[47135] == 47135 && 
b[47136] == 47136 && 
b[47137] == 47137 && 
b[47138] == 47138 && 
b[47139] == 47139 && 
b[47140] == 47140 && 
b[47141] == 47141 && 
b[47142] == 47142 && 
b[47143] == 47143 && 
b[47144] == 47144 && 
b[47145] == 47145 && 
b[47146] == 47146 && 
b[47147] == 47147 && 
b[47148] == 47148 && 
b[47149] == 47149 && 
b[47150] == 47150 && 
b[47151] == 47151 && 
b[47152] == 47152 && 
b[47153] == 47153 && 
b[47154] == 47154 && 
b[47155] == 47155 && 
b[47156] == 47156 && 
b[47157] == 47157 && 
b[47158] == 47158 && 
b[47159] == 47159 && 
b[47160] == 47160 && 
b[47161] == 47161 && 
b[47162] == 47162 && 
b[47163] == 47163 && 
b[47164] == 47164 && 
b[47165] == 47165 && 
b[47166] == 47166 && 
b[47167] == 47167 && 
b[47168] == 47168 && 
b[47169] == 47169 && 
b[47170] == 47170 && 
b[47171] == 47171 && 
b[47172] == 47172 && 
b[47173] == 47173 && 
b[47174] == 47174 && 
b[47175] == 47175 && 
b[47176] == 47176 && 
b[47177] == 47177 && 
b[47178] == 47178 && 
b[47179] == 47179 && 
b[47180] == 47180 && 
b[47181] == 47181 && 
b[47182] == 47182 && 
b[47183] == 47183 && 
b[47184] == 47184 && 
b[47185] == 47185 && 
b[47186] == 47186 && 
b[47187] == 47187 && 
b[47188] == 47188 && 
b[47189] == 47189 && 
b[47190] == 47190 && 
b[47191] == 47191 && 
b[47192] == 47192 && 
b[47193] == 47193 && 
b[47194] == 47194 && 
b[47195] == 47195 && 
b[47196] == 47196 && 
b[47197] == 47197 && 
b[47198] == 47198 && 
b[47199] == 47199 && 
b[47200] == 47200 && 
b[47201] == 47201 && 
b[47202] == 47202 && 
b[47203] == 47203 && 
b[47204] == 47204 && 
b[47205] == 47205 && 
b[47206] == 47206 && 
b[47207] == 47207 && 
b[47208] == 47208 && 
b[47209] == 47209 && 
b[47210] == 47210 && 
b[47211] == 47211 && 
b[47212] == 47212 && 
b[47213] == 47213 && 
b[47214] == 47214 && 
b[47215] == 47215 && 
b[47216] == 47216 && 
b[47217] == 47217 && 
b[47218] == 47218 && 
b[47219] == 47219 && 
b[47220] == 47220 && 
b[47221] == 47221 && 
b[47222] == 47222 && 
b[47223] == 47223 && 
b[47224] == 47224 && 
b[47225] == 47225 && 
b[47226] == 47226 && 
b[47227] == 47227 && 
b[47228] == 47228 && 
b[47229] == 47229 && 
b[47230] == 47230 && 
b[47231] == 47231 && 
b[47232] == 47232 && 
b[47233] == 47233 && 
b[47234] == 47234 && 
b[47235] == 47235 && 
b[47236] == 47236 && 
b[47237] == 47237 && 
b[47238] == 47238 && 
b[47239] == 47239 && 
b[47240] == 47240 && 
b[47241] == 47241 && 
b[47242] == 47242 && 
b[47243] == 47243 && 
b[47244] == 47244 && 
b[47245] == 47245 && 
b[47246] == 47246 && 
b[47247] == 47247 && 
b[47248] == 47248 && 
b[47249] == 47249 && 
b[47250] == 47250 && 
b[47251] == 47251 && 
b[47252] == 47252 && 
b[47253] == 47253 && 
b[47254] == 47254 && 
b[47255] == 47255 && 
b[47256] == 47256 && 
b[47257] == 47257 && 
b[47258] == 47258 && 
b[47259] == 47259 && 
b[47260] == 47260 && 
b[47261] == 47261 && 
b[47262] == 47262 && 
b[47263] == 47263 && 
b[47264] == 47264 && 
b[47265] == 47265 && 
b[47266] == 47266 && 
b[47267] == 47267 && 
b[47268] == 47268 && 
b[47269] == 47269 && 
b[47270] == 47270 && 
b[47271] == 47271 && 
b[47272] == 47272 && 
b[47273] == 47273 && 
b[47274] == 47274 && 
b[47275] == 47275 && 
b[47276] == 47276 && 
b[47277] == 47277 && 
b[47278] == 47278 && 
b[47279] == 47279 && 
b[47280] == 47280 && 
b[47281] == 47281 && 
b[47282] == 47282 && 
b[47283] == 47283 && 
b[47284] == 47284 && 
b[47285] == 47285 && 
b[47286] == 47286 && 
b[47287] == 47287 && 
b[47288] == 47288 && 
b[47289] == 47289 && 
b[47290] == 47290 && 
b[47291] == 47291 && 
b[47292] == 47292 && 
b[47293] == 47293 && 
b[47294] == 47294 && 
b[47295] == 47295 && 
b[47296] == 47296 && 
b[47297] == 47297 && 
b[47298] == 47298 && 
b[47299] == 47299 && 
b[47300] == 47300 && 
b[47301] == 47301 && 
b[47302] == 47302 && 
b[47303] == 47303 && 
b[47304] == 47304 && 
b[47305] == 47305 && 
b[47306] == 47306 && 
b[47307] == 47307 && 
b[47308] == 47308 && 
b[47309] == 47309 && 
b[47310] == 47310 && 
b[47311] == 47311 && 
b[47312] == 47312 && 
b[47313] == 47313 && 
b[47314] == 47314 && 
b[47315] == 47315 && 
b[47316] == 47316 && 
b[47317] == 47317 && 
b[47318] == 47318 && 
b[47319] == 47319 && 
b[47320] == 47320 && 
b[47321] == 47321 && 
b[47322] == 47322 && 
b[47323] == 47323 && 
b[47324] == 47324 && 
b[47325] == 47325 && 
b[47326] == 47326 && 
b[47327] == 47327 && 
b[47328] == 47328 && 
b[47329] == 47329 && 
b[47330] == 47330 && 
b[47331] == 47331 && 
b[47332] == 47332 && 
b[47333] == 47333 && 
b[47334] == 47334 && 
b[47335] == 47335 && 
b[47336] == 47336 && 
b[47337] == 47337 && 
b[47338] == 47338 && 
b[47339] == 47339 && 
b[47340] == 47340 && 
b[47341] == 47341 && 
b[47342] == 47342 && 
b[47343] == 47343 && 
b[47344] == 47344 && 
b[47345] == 47345 && 
b[47346] == 47346 && 
b[47347] == 47347 && 
b[47348] == 47348 && 
b[47349] == 47349 && 
b[47350] == 47350 && 
b[47351] == 47351 && 
b[47352] == 47352 && 
b[47353] == 47353 && 
b[47354] == 47354 && 
b[47355] == 47355 && 
b[47356] == 47356 && 
b[47357] == 47357 && 
b[47358] == 47358 && 
b[47359] == 47359 && 
b[47360] == 47360 && 
b[47361] == 47361 && 
b[47362] == 47362 && 
b[47363] == 47363 && 
b[47364] == 47364 && 
b[47365] == 47365 && 
b[47366] == 47366 && 
b[47367] == 47367 && 
b[47368] == 47368 && 
b[47369] == 47369 && 
b[47370] == 47370 && 
b[47371] == 47371 && 
b[47372] == 47372 && 
b[47373] == 47373 && 
b[47374] == 47374 && 
b[47375] == 47375 && 
b[47376] == 47376 && 
b[47377] == 47377 && 
b[47378] == 47378 && 
b[47379] == 47379 && 
b[47380] == 47380 && 
b[47381] == 47381 && 
b[47382] == 47382 && 
b[47383] == 47383 && 
b[47384] == 47384 && 
b[47385] == 47385 && 
b[47386] == 47386 && 
b[47387] == 47387 && 
b[47388] == 47388 && 
b[47389] == 47389 && 
b[47390] == 47390 && 
b[47391] == 47391 && 
b[47392] == 47392 && 
b[47393] == 47393 && 
b[47394] == 47394 && 
b[47395] == 47395 && 
b[47396] == 47396 && 
b[47397] == 47397 && 
b[47398] == 47398 && 
b[47399] == 47399 && 
b[47400] == 47400 && 
b[47401] == 47401 && 
b[47402] == 47402 && 
b[47403] == 47403 && 
b[47404] == 47404 && 
b[47405] == 47405 && 
b[47406] == 47406 && 
b[47407] == 47407 && 
b[47408] == 47408 && 
b[47409] == 47409 && 
b[47410] == 47410 && 
b[47411] == 47411 && 
b[47412] == 47412 && 
b[47413] == 47413 && 
b[47414] == 47414 && 
b[47415] == 47415 && 
b[47416] == 47416 && 
b[47417] == 47417 && 
b[47418] == 47418 && 
b[47419] == 47419 && 
b[47420] == 47420 && 
b[47421] == 47421 && 
b[47422] == 47422 && 
b[47423] == 47423 && 
b[47424] == 47424 && 
b[47425] == 47425 && 
b[47426] == 47426 && 
b[47427] == 47427 && 
b[47428] == 47428 && 
b[47429] == 47429 && 
b[47430] == 47430 && 
b[47431] == 47431 && 
b[47432] == 47432 && 
b[47433] == 47433 && 
b[47434] == 47434 && 
b[47435] == 47435 && 
b[47436] == 47436 && 
b[47437] == 47437 && 
b[47438] == 47438 && 
b[47439] == 47439 && 
b[47440] == 47440 && 
b[47441] == 47441 && 
b[47442] == 47442 && 
b[47443] == 47443 && 
b[47444] == 47444 && 
b[47445] == 47445 && 
b[47446] == 47446 && 
b[47447] == 47447 && 
b[47448] == 47448 && 
b[47449] == 47449 && 
b[47450] == 47450 && 
b[47451] == 47451 && 
b[47452] == 47452 && 
b[47453] == 47453 && 
b[47454] == 47454 && 
b[47455] == 47455 && 
b[47456] == 47456 && 
b[47457] == 47457 && 
b[47458] == 47458 && 
b[47459] == 47459 && 
b[47460] == 47460 && 
b[47461] == 47461 && 
b[47462] == 47462 && 
b[47463] == 47463 && 
b[47464] == 47464 && 
b[47465] == 47465 && 
b[47466] == 47466 && 
b[47467] == 47467 && 
b[47468] == 47468 && 
b[47469] == 47469 && 
b[47470] == 47470 && 
b[47471] == 47471 && 
b[47472] == 47472 && 
b[47473] == 47473 && 
b[47474] == 47474 && 
b[47475] == 47475 && 
b[47476] == 47476 && 
b[47477] == 47477 && 
b[47478] == 47478 && 
b[47479] == 47479 && 
b[47480] == 47480 && 
b[47481] == 47481 && 
b[47482] == 47482 && 
b[47483] == 47483 && 
b[47484] == 47484 && 
b[47485] == 47485 && 
b[47486] == 47486 && 
b[47487] == 47487 && 
b[47488] == 47488 && 
b[47489] == 47489 && 
b[47490] == 47490 && 
b[47491] == 47491 && 
b[47492] == 47492 && 
b[47493] == 47493 && 
b[47494] == 47494 && 
b[47495] == 47495 && 
b[47496] == 47496 && 
b[47497] == 47497 && 
b[47498] == 47498 && 
b[47499] == 47499 && 
b[47500] == 47500 && 
b[47501] == 47501 && 
b[47502] == 47502 && 
b[47503] == 47503 && 
b[47504] == 47504 && 
b[47505] == 47505 && 
b[47506] == 47506 && 
b[47507] == 47507 && 
b[47508] == 47508 && 
b[47509] == 47509 && 
b[47510] == 47510 && 
b[47511] == 47511 && 
b[47512] == 47512 && 
b[47513] == 47513 && 
b[47514] == 47514 && 
b[47515] == 47515 && 
b[47516] == 47516 && 
b[47517] == 47517 && 
b[47518] == 47518 && 
b[47519] == 47519 && 
b[47520] == 47520 && 
b[47521] == 47521 && 
b[47522] == 47522 && 
b[47523] == 47523 && 
b[47524] == 47524 && 
b[47525] == 47525 && 
b[47526] == 47526 && 
b[47527] == 47527 && 
b[47528] == 47528 && 
b[47529] == 47529 && 
b[47530] == 47530 && 
b[47531] == 47531 && 
b[47532] == 47532 && 
b[47533] == 47533 && 
b[47534] == 47534 && 
b[47535] == 47535 && 
b[47536] == 47536 && 
b[47537] == 47537 && 
b[47538] == 47538 && 
b[47539] == 47539 && 
b[47540] == 47540 && 
b[47541] == 47541 && 
b[47542] == 47542 && 
b[47543] == 47543 && 
b[47544] == 47544 && 
b[47545] == 47545 && 
b[47546] == 47546 && 
b[47547] == 47547 && 
b[47548] == 47548 && 
b[47549] == 47549 && 
b[47550] == 47550 && 
b[47551] == 47551 && 
b[47552] == 47552 && 
b[47553] == 47553 && 
b[47554] == 47554 && 
b[47555] == 47555 && 
b[47556] == 47556 && 
b[47557] == 47557 && 
b[47558] == 47558 && 
b[47559] == 47559 && 
b[47560] == 47560 && 
b[47561] == 47561 && 
b[47562] == 47562 && 
b[47563] == 47563 && 
b[47564] == 47564 && 
b[47565] == 47565 && 
b[47566] == 47566 && 
b[47567] == 47567 && 
b[47568] == 47568 && 
b[47569] == 47569 && 
b[47570] == 47570 && 
b[47571] == 47571 && 
b[47572] == 47572 && 
b[47573] == 47573 && 
b[47574] == 47574 && 
b[47575] == 47575 && 
b[47576] == 47576 && 
b[47577] == 47577 && 
b[47578] == 47578 && 
b[47579] == 47579 && 
b[47580] == 47580 && 
b[47581] == 47581 && 
b[47582] == 47582 && 
b[47583] == 47583 && 
b[47584] == 47584 && 
b[47585] == 47585 && 
b[47586] == 47586 && 
b[47587] == 47587 && 
b[47588] == 47588 && 
b[47589] == 47589 && 
b[47590] == 47590 && 
b[47591] == 47591 && 
b[47592] == 47592 && 
b[47593] == 47593 && 
b[47594] == 47594 && 
b[47595] == 47595 && 
b[47596] == 47596 && 
b[47597] == 47597 && 
b[47598] == 47598 && 
b[47599] == 47599 && 
b[47600] == 47600 && 
b[47601] == 47601 && 
b[47602] == 47602 && 
b[47603] == 47603 && 
b[47604] == 47604 && 
b[47605] == 47605 && 
b[47606] == 47606 && 
b[47607] == 47607 && 
b[47608] == 47608 && 
b[47609] == 47609 && 
b[47610] == 47610 && 
b[47611] == 47611 && 
b[47612] == 47612 && 
b[47613] == 47613 && 
b[47614] == 47614 && 
b[47615] == 47615 && 
b[47616] == 47616 && 
b[47617] == 47617 && 
b[47618] == 47618 && 
b[47619] == 47619 && 
b[47620] == 47620 && 
b[47621] == 47621 && 
b[47622] == 47622 && 
b[47623] == 47623 && 
b[47624] == 47624 && 
b[47625] == 47625 && 
b[47626] == 47626 && 
b[47627] == 47627 && 
b[47628] == 47628 && 
b[47629] == 47629 && 
b[47630] == 47630 && 
b[47631] == 47631 && 
b[47632] == 47632 && 
b[47633] == 47633 && 
b[47634] == 47634 && 
b[47635] == 47635 && 
b[47636] == 47636 && 
b[47637] == 47637 && 
b[47638] == 47638 && 
b[47639] == 47639 && 
b[47640] == 47640 && 
b[47641] == 47641 && 
b[47642] == 47642 && 
b[47643] == 47643 && 
b[47644] == 47644 && 
b[47645] == 47645 && 
b[47646] == 47646 && 
b[47647] == 47647 && 
b[47648] == 47648 && 
b[47649] == 47649 && 
b[47650] == 47650 && 
b[47651] == 47651 && 
b[47652] == 47652 && 
b[47653] == 47653 && 
b[47654] == 47654 && 
b[47655] == 47655 && 
b[47656] == 47656 && 
b[47657] == 47657 && 
b[47658] == 47658 && 
b[47659] == 47659 && 
b[47660] == 47660 && 
b[47661] == 47661 && 
b[47662] == 47662 && 
b[47663] == 47663 && 
b[47664] == 47664 && 
b[47665] == 47665 && 
b[47666] == 47666 && 
b[47667] == 47667 && 
b[47668] == 47668 && 
b[47669] == 47669 && 
b[47670] == 47670 && 
b[47671] == 47671 && 
b[47672] == 47672 && 
b[47673] == 47673 && 
b[47674] == 47674 && 
b[47675] == 47675 && 
b[47676] == 47676 && 
b[47677] == 47677 && 
b[47678] == 47678 && 
b[47679] == 47679 && 
b[47680] == 47680 && 
b[47681] == 47681 && 
b[47682] == 47682 && 
b[47683] == 47683 && 
b[47684] == 47684 && 
b[47685] == 47685 && 
b[47686] == 47686 && 
b[47687] == 47687 && 
b[47688] == 47688 && 
b[47689] == 47689 && 
b[47690] == 47690 && 
b[47691] == 47691 && 
b[47692] == 47692 && 
b[47693] == 47693 && 
b[47694] == 47694 && 
b[47695] == 47695 && 
b[47696] == 47696 && 
b[47697] == 47697 && 
b[47698] == 47698 && 
b[47699] == 47699 && 
b[47700] == 47700 && 
b[47701] == 47701 && 
b[47702] == 47702 && 
b[47703] == 47703 && 
b[47704] == 47704 && 
b[47705] == 47705 && 
b[47706] == 47706 && 
b[47707] == 47707 && 
b[47708] == 47708 && 
b[47709] == 47709 && 
b[47710] == 47710 && 
b[47711] == 47711 && 
b[47712] == 47712 && 
b[47713] == 47713 && 
b[47714] == 47714 && 
b[47715] == 47715 && 
b[47716] == 47716 && 
b[47717] == 47717 && 
b[47718] == 47718 && 
b[47719] == 47719 && 
b[47720] == 47720 && 
b[47721] == 47721 && 
b[47722] == 47722 && 
b[47723] == 47723 && 
b[47724] == 47724 && 
b[47725] == 47725 && 
b[47726] == 47726 && 
b[47727] == 47727 && 
b[47728] == 47728 && 
b[47729] == 47729 && 
b[47730] == 47730 && 
b[47731] == 47731 && 
b[47732] == 47732 && 
b[47733] == 47733 && 
b[47734] == 47734 && 
b[47735] == 47735 && 
b[47736] == 47736 && 
b[47737] == 47737 && 
b[47738] == 47738 && 
b[47739] == 47739 && 
b[47740] == 47740 && 
b[47741] == 47741 && 
b[47742] == 47742 && 
b[47743] == 47743 && 
b[47744] == 47744 && 
b[47745] == 47745 && 
b[47746] == 47746 && 
b[47747] == 47747 && 
b[47748] == 47748 && 
b[47749] == 47749 && 
b[47750] == 47750 && 
b[47751] == 47751 && 
b[47752] == 47752 && 
b[47753] == 47753 && 
b[47754] == 47754 && 
b[47755] == 47755 && 
b[47756] == 47756 && 
b[47757] == 47757 && 
b[47758] == 47758 && 
b[47759] == 47759 && 
b[47760] == 47760 && 
b[47761] == 47761 && 
b[47762] == 47762 && 
b[47763] == 47763 && 
b[47764] == 47764 && 
b[47765] == 47765 && 
b[47766] == 47766 && 
b[47767] == 47767 && 
b[47768] == 47768 && 
b[47769] == 47769 && 
b[47770] == 47770 && 
b[47771] == 47771 && 
b[47772] == 47772 && 
b[47773] == 47773 && 
b[47774] == 47774 && 
b[47775] == 47775 && 
b[47776] == 47776 && 
b[47777] == 47777 && 
b[47778] == 47778 && 
b[47779] == 47779 && 
b[47780] == 47780 && 
b[47781] == 47781 && 
b[47782] == 47782 && 
b[47783] == 47783 && 
b[47784] == 47784 && 
b[47785] == 47785 && 
b[47786] == 47786 && 
b[47787] == 47787 && 
b[47788] == 47788 && 
b[47789] == 47789 && 
b[47790] == 47790 && 
b[47791] == 47791 && 
b[47792] == 47792 && 
b[47793] == 47793 && 
b[47794] == 47794 && 
b[47795] == 47795 && 
b[47796] == 47796 && 
b[47797] == 47797 && 
b[47798] == 47798 && 
b[47799] == 47799 && 
b[47800] == 47800 && 
b[47801] == 47801 && 
b[47802] == 47802 && 
b[47803] == 47803 && 
b[47804] == 47804 && 
b[47805] == 47805 && 
b[47806] == 47806 && 
b[47807] == 47807 && 
b[47808] == 47808 && 
b[47809] == 47809 && 
b[47810] == 47810 && 
b[47811] == 47811 && 
b[47812] == 47812 && 
b[47813] == 47813 && 
b[47814] == 47814 && 
b[47815] == 47815 && 
b[47816] == 47816 && 
b[47817] == 47817 && 
b[47818] == 47818 && 
b[47819] == 47819 && 
b[47820] == 47820 && 
b[47821] == 47821 && 
b[47822] == 47822 && 
b[47823] == 47823 && 
b[47824] == 47824 && 
b[47825] == 47825 && 
b[47826] == 47826 && 
b[47827] == 47827 && 
b[47828] == 47828 && 
b[47829] == 47829 && 
b[47830] == 47830 && 
b[47831] == 47831 && 
b[47832] == 47832 && 
b[47833] == 47833 && 
b[47834] == 47834 && 
b[47835] == 47835 && 
b[47836] == 47836 && 
b[47837] == 47837 && 
b[47838] == 47838 && 
b[47839] == 47839 && 
b[47840] == 47840 && 
b[47841] == 47841 && 
b[47842] == 47842 && 
b[47843] == 47843 && 
b[47844] == 47844 && 
b[47845] == 47845 && 
b[47846] == 47846 && 
b[47847] == 47847 && 
b[47848] == 47848 && 
b[47849] == 47849 && 
b[47850] == 47850 && 
b[47851] == 47851 && 
b[47852] == 47852 && 
b[47853] == 47853 && 
b[47854] == 47854 && 
b[47855] == 47855 && 
b[47856] == 47856 && 
b[47857] == 47857 && 
b[47858] == 47858 && 
b[47859] == 47859 && 
b[47860] == 47860 && 
b[47861] == 47861 && 
b[47862] == 47862 && 
b[47863] == 47863 && 
b[47864] == 47864 && 
b[47865] == 47865 && 
b[47866] == 47866 && 
b[47867] == 47867 && 
b[47868] == 47868 && 
b[47869] == 47869 && 
b[47870] == 47870 && 
b[47871] == 47871 && 
b[47872] == 47872 && 
b[47873] == 47873 && 
b[47874] == 47874 && 
b[47875] == 47875 && 
b[47876] == 47876 && 
b[47877] == 47877 && 
b[47878] == 47878 && 
b[47879] == 47879 && 
b[47880] == 47880 && 
b[47881] == 47881 && 
b[47882] == 47882 && 
b[47883] == 47883 && 
b[47884] == 47884 && 
b[47885] == 47885 && 
b[47886] == 47886 && 
b[47887] == 47887 && 
b[47888] == 47888 && 
b[47889] == 47889 && 
b[47890] == 47890 && 
b[47891] == 47891 && 
b[47892] == 47892 && 
b[47893] == 47893 && 
b[47894] == 47894 && 
b[47895] == 47895 && 
b[47896] == 47896 && 
b[47897] == 47897 && 
b[47898] == 47898 && 
b[47899] == 47899 && 
b[47900] == 47900 && 
b[47901] == 47901 && 
b[47902] == 47902 && 
b[47903] == 47903 && 
b[47904] == 47904 && 
b[47905] == 47905 && 
b[47906] == 47906 && 
b[47907] == 47907 && 
b[47908] == 47908 && 
b[47909] == 47909 && 
b[47910] == 47910 && 
b[47911] == 47911 && 
b[47912] == 47912 && 
b[47913] == 47913 && 
b[47914] == 47914 && 
b[47915] == 47915 && 
b[47916] == 47916 && 
b[47917] == 47917 && 
b[47918] == 47918 && 
b[47919] == 47919 && 
b[47920] == 47920 && 
b[47921] == 47921 && 
b[47922] == 47922 && 
b[47923] == 47923 && 
b[47924] == 47924 && 
b[47925] == 47925 && 
b[47926] == 47926 && 
b[47927] == 47927 && 
b[47928] == 47928 && 
b[47929] == 47929 && 
b[47930] == 47930 && 
b[47931] == 47931 && 
b[47932] == 47932 && 
b[47933] == 47933 && 
b[47934] == 47934 && 
b[47935] == 47935 && 
b[47936] == 47936 && 
b[47937] == 47937 && 
b[47938] == 47938 && 
b[47939] == 47939 && 
b[47940] == 47940 && 
b[47941] == 47941 && 
b[47942] == 47942 && 
b[47943] == 47943 && 
b[47944] == 47944 && 
b[47945] == 47945 && 
b[47946] == 47946 && 
b[47947] == 47947 && 
b[47948] == 47948 && 
b[47949] == 47949 && 
b[47950] == 47950 && 
b[47951] == 47951 && 
b[47952] == 47952 && 
b[47953] == 47953 && 
b[47954] == 47954 && 
b[47955] == 47955 && 
b[47956] == 47956 && 
b[47957] == 47957 && 
b[47958] == 47958 && 
b[47959] == 47959 && 
b[47960] == 47960 && 
b[47961] == 47961 && 
b[47962] == 47962 && 
b[47963] == 47963 && 
b[47964] == 47964 && 
b[47965] == 47965 && 
b[47966] == 47966 && 
b[47967] == 47967 && 
b[47968] == 47968 && 
b[47969] == 47969 && 
b[47970] == 47970 && 
b[47971] == 47971 && 
b[47972] == 47972 && 
b[47973] == 47973 && 
b[47974] == 47974 && 
b[47975] == 47975 && 
b[47976] == 47976 && 
b[47977] == 47977 && 
b[47978] == 47978 && 
b[47979] == 47979 && 
b[47980] == 47980 && 
b[47981] == 47981 && 
b[47982] == 47982 && 
b[47983] == 47983 && 
b[47984] == 47984 && 
b[47985] == 47985 && 
b[47986] == 47986 && 
b[47987] == 47987 && 
b[47988] == 47988 && 
b[47989] == 47989 && 
b[47990] == 47990 && 
b[47991] == 47991 && 
b[47992] == 47992 && 
b[47993] == 47993 && 
b[47994] == 47994 && 
b[47995] == 47995 && 
b[47996] == 47996 && 
b[47997] == 47997 && 
b[47998] == 47998 && 
b[47999] == 47999 && 
b[48000] == 48000 && 
b[48001] == 48001 && 
b[48002] == 48002 && 
b[48003] == 48003 && 
b[48004] == 48004 && 
b[48005] == 48005 && 
b[48006] == 48006 && 
b[48007] == 48007 && 
b[48008] == 48008 && 
b[48009] == 48009 && 
b[48010] == 48010 && 
b[48011] == 48011 && 
b[48012] == 48012 && 
b[48013] == 48013 && 
b[48014] == 48014 && 
b[48015] == 48015 && 
b[48016] == 48016 && 
b[48017] == 48017 && 
b[48018] == 48018 && 
b[48019] == 48019 && 
b[48020] == 48020 && 
b[48021] == 48021 && 
b[48022] == 48022 && 
b[48023] == 48023 && 
b[48024] == 48024 && 
b[48025] == 48025 && 
b[48026] == 48026 && 
b[48027] == 48027 && 
b[48028] == 48028 && 
b[48029] == 48029 && 
b[48030] == 48030 && 
b[48031] == 48031 && 
b[48032] == 48032 && 
b[48033] == 48033 && 
b[48034] == 48034 && 
b[48035] == 48035 && 
b[48036] == 48036 && 
b[48037] == 48037 && 
b[48038] == 48038 && 
b[48039] == 48039 && 
b[48040] == 48040 && 
b[48041] == 48041 && 
b[48042] == 48042 && 
b[48043] == 48043 && 
b[48044] == 48044 && 
b[48045] == 48045 && 
b[48046] == 48046 && 
b[48047] == 48047 && 
b[48048] == 48048 && 
b[48049] == 48049 && 
b[48050] == 48050 && 
b[48051] == 48051 && 
b[48052] == 48052 && 
b[48053] == 48053 && 
b[48054] == 48054 && 
b[48055] == 48055 && 
b[48056] == 48056 && 
b[48057] == 48057 && 
b[48058] == 48058 && 
b[48059] == 48059 && 
b[48060] == 48060 && 
b[48061] == 48061 && 
b[48062] == 48062 && 
b[48063] == 48063 && 
b[48064] == 48064 && 
b[48065] == 48065 && 
b[48066] == 48066 && 
b[48067] == 48067 && 
b[48068] == 48068 && 
b[48069] == 48069 && 
b[48070] == 48070 && 
b[48071] == 48071 && 
b[48072] == 48072 && 
b[48073] == 48073 && 
b[48074] == 48074 && 
b[48075] == 48075 && 
b[48076] == 48076 && 
b[48077] == 48077 && 
b[48078] == 48078 && 
b[48079] == 48079 && 
b[48080] == 48080 && 
b[48081] == 48081 && 
b[48082] == 48082 && 
b[48083] == 48083 && 
b[48084] == 48084 && 
b[48085] == 48085 && 
b[48086] == 48086 && 
b[48087] == 48087 && 
b[48088] == 48088 && 
b[48089] == 48089 && 
b[48090] == 48090 && 
b[48091] == 48091 && 
b[48092] == 48092 && 
b[48093] == 48093 && 
b[48094] == 48094 && 
b[48095] == 48095 && 
b[48096] == 48096 && 
b[48097] == 48097 && 
b[48098] == 48098 && 
b[48099] == 48099 && 
b[48100] == 48100 && 
b[48101] == 48101 && 
b[48102] == 48102 && 
b[48103] == 48103 && 
b[48104] == 48104 && 
b[48105] == 48105 && 
b[48106] == 48106 && 
b[48107] == 48107 && 
b[48108] == 48108 && 
b[48109] == 48109 && 
b[48110] == 48110 && 
b[48111] == 48111 && 
b[48112] == 48112 && 
b[48113] == 48113 && 
b[48114] == 48114 && 
b[48115] == 48115 && 
b[48116] == 48116 && 
b[48117] == 48117 && 
b[48118] == 48118 && 
b[48119] == 48119 && 
b[48120] == 48120 && 
b[48121] == 48121 && 
b[48122] == 48122 && 
b[48123] == 48123 && 
b[48124] == 48124 && 
b[48125] == 48125 && 
b[48126] == 48126 && 
b[48127] == 48127 && 
b[48128] == 48128 && 
b[48129] == 48129 && 
b[48130] == 48130 && 
b[48131] == 48131 && 
b[48132] == 48132 && 
b[48133] == 48133 && 
b[48134] == 48134 && 
b[48135] == 48135 && 
b[48136] == 48136 && 
b[48137] == 48137 && 
b[48138] == 48138 && 
b[48139] == 48139 && 
b[48140] == 48140 && 
b[48141] == 48141 && 
b[48142] == 48142 && 
b[48143] == 48143 && 
b[48144] == 48144 && 
b[48145] == 48145 && 
b[48146] == 48146 && 
b[48147] == 48147 && 
b[48148] == 48148 && 
b[48149] == 48149 && 
b[48150] == 48150 && 
b[48151] == 48151 && 
b[48152] == 48152 && 
b[48153] == 48153 && 
b[48154] == 48154 && 
b[48155] == 48155 && 
b[48156] == 48156 && 
b[48157] == 48157 && 
b[48158] == 48158 && 
b[48159] == 48159 && 
b[48160] == 48160 && 
b[48161] == 48161 && 
b[48162] == 48162 && 
b[48163] == 48163 && 
b[48164] == 48164 && 
b[48165] == 48165 && 
b[48166] == 48166 && 
b[48167] == 48167 && 
b[48168] == 48168 && 
b[48169] == 48169 && 
b[48170] == 48170 && 
b[48171] == 48171 && 
b[48172] == 48172 && 
b[48173] == 48173 && 
b[48174] == 48174 && 
b[48175] == 48175 && 
b[48176] == 48176 && 
b[48177] == 48177 && 
b[48178] == 48178 && 
b[48179] == 48179 && 
b[48180] == 48180 && 
b[48181] == 48181 && 
b[48182] == 48182 && 
b[48183] == 48183 && 
b[48184] == 48184 && 
b[48185] == 48185 && 
b[48186] == 48186 && 
b[48187] == 48187 && 
b[48188] == 48188 && 
b[48189] == 48189 && 
b[48190] == 48190 && 
b[48191] == 48191 && 
b[48192] == 48192 && 
b[48193] == 48193 && 
b[48194] == 48194 && 
b[48195] == 48195 && 
b[48196] == 48196 && 
b[48197] == 48197 && 
b[48198] == 48198 && 
b[48199] == 48199 && 
b[48200] == 48200 && 
b[48201] == 48201 && 
b[48202] == 48202 && 
b[48203] == 48203 && 
b[48204] == 48204 && 
b[48205] == 48205 && 
b[48206] == 48206 && 
b[48207] == 48207 && 
b[48208] == 48208 && 
b[48209] == 48209 && 
b[48210] == 48210 && 
b[48211] == 48211 && 
b[48212] == 48212 && 
b[48213] == 48213 && 
b[48214] == 48214 && 
b[48215] == 48215 && 
b[48216] == 48216 && 
b[48217] == 48217 && 
b[48218] == 48218 && 
b[48219] == 48219 && 
b[48220] == 48220 && 
b[48221] == 48221 && 
b[48222] == 48222 && 
b[48223] == 48223 && 
b[48224] == 48224 && 
b[48225] == 48225 && 
b[48226] == 48226 && 
b[48227] == 48227 && 
b[48228] == 48228 && 
b[48229] == 48229 && 
b[48230] == 48230 && 
b[48231] == 48231 && 
b[48232] == 48232 && 
b[48233] == 48233 && 
b[48234] == 48234 && 
b[48235] == 48235 && 
b[48236] == 48236 && 
b[48237] == 48237 && 
b[48238] == 48238 && 
b[48239] == 48239 && 
b[48240] == 48240 && 
b[48241] == 48241 && 
b[48242] == 48242 && 
b[48243] == 48243 && 
b[48244] == 48244 && 
b[48245] == 48245 && 
b[48246] == 48246 && 
b[48247] == 48247 && 
b[48248] == 48248 && 
b[48249] == 48249 && 
b[48250] == 48250 && 
b[48251] == 48251 && 
b[48252] == 48252 && 
b[48253] == 48253 && 
b[48254] == 48254 && 
b[48255] == 48255 && 
b[48256] == 48256 && 
b[48257] == 48257 && 
b[48258] == 48258 && 
b[48259] == 48259 && 
b[48260] == 48260 && 
b[48261] == 48261 && 
b[48262] == 48262 && 
b[48263] == 48263 && 
b[48264] == 48264 && 
b[48265] == 48265 && 
b[48266] == 48266 && 
b[48267] == 48267 && 
b[48268] == 48268 && 
b[48269] == 48269 && 
b[48270] == 48270 && 
b[48271] == 48271 && 
b[48272] == 48272 && 
b[48273] == 48273 && 
b[48274] == 48274 && 
b[48275] == 48275 && 
b[48276] == 48276 && 
b[48277] == 48277 && 
b[48278] == 48278 && 
b[48279] == 48279 && 
b[48280] == 48280 && 
b[48281] == 48281 && 
b[48282] == 48282 && 
b[48283] == 48283 && 
b[48284] == 48284 && 
b[48285] == 48285 && 
b[48286] == 48286 && 
b[48287] == 48287 && 
b[48288] == 48288 && 
b[48289] == 48289 && 
b[48290] == 48290 && 
b[48291] == 48291 && 
b[48292] == 48292 && 
b[48293] == 48293 && 
b[48294] == 48294 && 
b[48295] == 48295 && 
b[48296] == 48296 && 
b[48297] == 48297 && 
b[48298] == 48298 && 
b[48299] == 48299 && 
b[48300] == 48300 && 
b[48301] == 48301 && 
b[48302] == 48302 && 
b[48303] == 48303 && 
b[48304] == 48304 && 
b[48305] == 48305 && 
b[48306] == 48306 && 
b[48307] == 48307 && 
b[48308] == 48308 && 
b[48309] == 48309 && 
b[48310] == 48310 && 
b[48311] == 48311 && 
b[48312] == 48312 && 
b[48313] == 48313 && 
b[48314] == 48314 && 
b[48315] == 48315 && 
b[48316] == 48316 && 
b[48317] == 48317 && 
b[48318] == 48318 && 
b[48319] == 48319 && 
b[48320] == 48320 && 
b[48321] == 48321 && 
b[48322] == 48322 && 
b[48323] == 48323 && 
b[48324] == 48324 && 
b[48325] == 48325 && 
b[48326] == 48326 && 
b[48327] == 48327 && 
b[48328] == 48328 && 
b[48329] == 48329 && 
b[48330] == 48330 && 
b[48331] == 48331 && 
b[48332] == 48332 && 
b[48333] == 48333 && 
b[48334] == 48334 && 
b[48335] == 48335 && 
b[48336] == 48336 && 
b[48337] == 48337 && 
b[48338] == 48338 && 
b[48339] == 48339 && 
b[48340] == 48340 && 
b[48341] == 48341 && 
b[48342] == 48342 && 
b[48343] == 48343 && 
b[48344] == 48344 && 
b[48345] == 48345 && 
b[48346] == 48346 && 
b[48347] == 48347 && 
b[48348] == 48348 && 
b[48349] == 48349 && 
b[48350] == 48350 && 
b[48351] == 48351 && 
b[48352] == 48352 && 
b[48353] == 48353 && 
b[48354] == 48354 && 
b[48355] == 48355 && 
b[48356] == 48356 && 
b[48357] == 48357 && 
b[48358] == 48358 && 
b[48359] == 48359 && 
b[48360] == 48360 && 
b[48361] == 48361 && 
b[48362] == 48362 && 
b[48363] == 48363 && 
b[48364] == 48364 && 
b[48365] == 48365 && 
b[48366] == 48366 && 
b[48367] == 48367 && 
b[48368] == 48368 && 
b[48369] == 48369 && 
b[48370] == 48370 && 
b[48371] == 48371 && 
b[48372] == 48372 && 
b[48373] == 48373 && 
b[48374] == 48374 && 
b[48375] == 48375 && 
b[48376] == 48376 && 
b[48377] == 48377 && 
b[48378] == 48378 && 
b[48379] == 48379 && 
b[48380] == 48380 && 
b[48381] == 48381 && 
b[48382] == 48382 && 
b[48383] == 48383 && 
b[48384] == 48384 && 
b[48385] == 48385 && 
b[48386] == 48386 && 
b[48387] == 48387 && 
b[48388] == 48388 && 
b[48389] == 48389 && 
b[48390] == 48390 && 
b[48391] == 48391 && 
b[48392] == 48392 && 
b[48393] == 48393 && 
b[48394] == 48394 && 
b[48395] == 48395 && 
b[48396] == 48396 && 
b[48397] == 48397 && 
b[48398] == 48398 && 
b[48399] == 48399 && 
b[48400] == 48400 && 
b[48401] == 48401 && 
b[48402] == 48402 && 
b[48403] == 48403 && 
b[48404] == 48404 && 
b[48405] == 48405 && 
b[48406] == 48406 && 
b[48407] == 48407 && 
b[48408] == 48408 && 
b[48409] == 48409 && 
b[48410] == 48410 && 
b[48411] == 48411 && 
b[48412] == 48412 && 
b[48413] == 48413 && 
b[48414] == 48414 && 
b[48415] == 48415 && 
b[48416] == 48416 && 
b[48417] == 48417 && 
b[48418] == 48418 && 
b[48419] == 48419 && 
b[48420] == 48420 && 
b[48421] == 48421 && 
b[48422] == 48422 && 
b[48423] == 48423 && 
b[48424] == 48424 && 
b[48425] == 48425 && 
b[48426] == 48426 && 
b[48427] == 48427 && 
b[48428] == 48428 && 
b[48429] == 48429 && 
b[48430] == 48430 && 
b[48431] == 48431 && 
b[48432] == 48432 && 
b[48433] == 48433 && 
b[48434] == 48434 && 
b[48435] == 48435 && 
b[48436] == 48436 && 
b[48437] == 48437 && 
b[48438] == 48438 && 
b[48439] == 48439 && 
b[48440] == 48440 && 
b[48441] == 48441 && 
b[48442] == 48442 && 
b[48443] == 48443 && 
b[48444] == 48444 && 
b[48445] == 48445 && 
b[48446] == 48446 && 
b[48447] == 48447 && 
b[48448] == 48448 && 
b[48449] == 48449 && 
b[48450] == 48450 && 
b[48451] == 48451 && 
b[48452] == 48452 && 
b[48453] == 48453 && 
b[48454] == 48454 && 
b[48455] == 48455 && 
b[48456] == 48456 && 
b[48457] == 48457 && 
b[48458] == 48458 && 
b[48459] == 48459 && 
b[48460] == 48460 && 
b[48461] == 48461 && 
b[48462] == 48462 && 
b[48463] == 48463 && 
b[48464] == 48464 && 
b[48465] == 48465 && 
b[48466] == 48466 && 
b[48467] == 48467 && 
b[48468] == 48468 && 
b[48469] == 48469 && 
b[48470] == 48470 && 
b[48471] == 48471 && 
b[48472] == 48472 && 
b[48473] == 48473 && 
b[48474] == 48474 && 
b[48475] == 48475 && 
b[48476] == 48476 && 
b[48477] == 48477 && 
b[48478] == 48478 && 
b[48479] == 48479 && 
b[48480] == 48480 && 
b[48481] == 48481 && 
b[48482] == 48482 && 
b[48483] == 48483 && 
b[48484] == 48484 && 
b[48485] == 48485 && 
b[48486] == 48486 && 
b[48487] == 48487 && 
b[48488] == 48488 && 
b[48489] == 48489 && 
b[48490] == 48490 && 
b[48491] == 48491 && 
b[48492] == 48492 && 
b[48493] == 48493 && 
b[48494] == 48494 && 
b[48495] == 48495 && 
b[48496] == 48496 && 
b[48497] == 48497 && 
b[48498] == 48498 && 
b[48499] == 48499 && 
b[48500] == 48500 && 
b[48501] == 48501 && 
b[48502] == 48502 && 
b[48503] == 48503 && 
b[48504] == 48504 && 
b[48505] == 48505 && 
b[48506] == 48506 && 
b[48507] == 48507 && 
b[48508] == 48508 && 
b[48509] == 48509 && 
b[48510] == 48510 && 
b[48511] == 48511 && 
b[48512] == 48512 && 
b[48513] == 48513 && 
b[48514] == 48514 && 
b[48515] == 48515 && 
b[48516] == 48516 && 
b[48517] == 48517 && 
b[48518] == 48518 && 
b[48519] == 48519 && 
b[48520] == 48520 && 
b[48521] == 48521 && 
b[48522] == 48522 && 
b[48523] == 48523 && 
b[48524] == 48524 && 
b[48525] == 48525 && 
b[48526] == 48526 && 
b[48527] == 48527 && 
b[48528] == 48528 && 
b[48529] == 48529 && 
b[48530] == 48530 && 
b[48531] == 48531 && 
b[48532] == 48532 && 
b[48533] == 48533 && 
b[48534] == 48534 && 
b[48535] == 48535 && 
b[48536] == 48536 && 
b[48537] == 48537 && 
b[48538] == 48538 && 
b[48539] == 48539 && 
b[48540] == 48540 && 
b[48541] == 48541 && 
b[48542] == 48542 && 
b[48543] == 48543 && 
b[48544] == 48544 && 
b[48545] == 48545 && 
b[48546] == 48546 && 
b[48547] == 48547 && 
b[48548] == 48548 && 
b[48549] == 48549 && 
b[48550] == 48550 && 
b[48551] == 48551 && 
b[48552] == 48552 && 
b[48553] == 48553 && 
b[48554] == 48554 && 
b[48555] == 48555 && 
b[48556] == 48556 && 
b[48557] == 48557 && 
b[48558] == 48558 && 
b[48559] == 48559 && 
b[48560] == 48560 && 
b[48561] == 48561 && 
b[48562] == 48562 && 
b[48563] == 48563 && 
b[48564] == 48564 && 
b[48565] == 48565 && 
b[48566] == 48566 && 
b[48567] == 48567 && 
b[48568] == 48568 && 
b[48569] == 48569 && 
b[48570] == 48570 && 
b[48571] == 48571 && 
b[48572] == 48572 && 
b[48573] == 48573 && 
b[48574] == 48574 && 
b[48575] == 48575 && 
b[48576] == 48576 && 
b[48577] == 48577 && 
b[48578] == 48578 && 
b[48579] == 48579 && 
b[48580] == 48580 && 
b[48581] == 48581 && 
b[48582] == 48582 && 
b[48583] == 48583 && 
b[48584] == 48584 && 
b[48585] == 48585 && 
b[48586] == 48586 && 
b[48587] == 48587 && 
b[48588] == 48588 && 
b[48589] == 48589 && 
b[48590] == 48590 && 
b[48591] == 48591 && 
b[48592] == 48592 && 
b[48593] == 48593 && 
b[48594] == 48594 && 
b[48595] == 48595 && 
b[48596] == 48596 && 
b[48597] == 48597 && 
b[48598] == 48598 && 
b[48599] == 48599 && 
b[48600] == 48600 && 
b[48601] == 48601 && 
b[48602] == 48602 && 
b[48603] == 48603 && 
b[48604] == 48604 && 
b[48605] == 48605 && 
b[48606] == 48606 && 
b[48607] == 48607 && 
b[48608] == 48608 && 
b[48609] == 48609 && 
b[48610] == 48610 && 
b[48611] == 48611 && 
b[48612] == 48612 && 
b[48613] == 48613 && 
b[48614] == 48614 && 
b[48615] == 48615 && 
b[48616] == 48616 && 
b[48617] == 48617 && 
b[48618] == 48618 && 
b[48619] == 48619 && 
b[48620] == 48620 && 
b[48621] == 48621 && 
b[48622] == 48622 && 
b[48623] == 48623 && 
b[48624] == 48624 && 
b[48625] == 48625 && 
b[48626] == 48626 && 
b[48627] == 48627 && 
b[48628] == 48628 && 
b[48629] == 48629 && 
b[48630] == 48630 && 
b[48631] == 48631 && 
b[48632] == 48632 && 
b[48633] == 48633 && 
b[48634] == 48634 && 
b[48635] == 48635 && 
b[48636] == 48636 && 
b[48637] == 48637 && 
b[48638] == 48638 && 
b[48639] == 48639 && 
b[48640] == 48640 && 
b[48641] == 48641 && 
b[48642] == 48642 && 
b[48643] == 48643 && 
b[48644] == 48644 && 
b[48645] == 48645 && 
b[48646] == 48646 && 
b[48647] == 48647 && 
b[48648] == 48648 && 
b[48649] == 48649 && 
b[48650] == 48650 && 
b[48651] == 48651 && 
b[48652] == 48652 && 
b[48653] == 48653 && 
b[48654] == 48654 && 
b[48655] == 48655 && 
b[48656] == 48656 && 
b[48657] == 48657 && 
b[48658] == 48658 && 
b[48659] == 48659 && 
b[48660] == 48660 && 
b[48661] == 48661 && 
b[48662] == 48662 && 
b[48663] == 48663 && 
b[48664] == 48664 && 
b[48665] == 48665 && 
b[48666] == 48666 && 
b[48667] == 48667 && 
b[48668] == 48668 && 
b[48669] == 48669 && 
b[48670] == 48670 && 
b[48671] == 48671 && 
b[48672] == 48672 && 
b[48673] == 48673 && 
b[48674] == 48674 && 
b[48675] == 48675 && 
b[48676] == 48676 && 
b[48677] == 48677 && 
b[48678] == 48678 && 
b[48679] == 48679 && 
b[48680] == 48680 && 
b[48681] == 48681 && 
b[48682] == 48682 && 
b[48683] == 48683 && 
b[48684] == 48684 && 
b[48685] == 48685 && 
b[48686] == 48686 && 
b[48687] == 48687 && 
b[48688] == 48688 && 
b[48689] == 48689 && 
b[48690] == 48690 && 
b[48691] == 48691 && 
b[48692] == 48692 && 
b[48693] == 48693 && 
b[48694] == 48694 && 
b[48695] == 48695 && 
b[48696] == 48696 && 
b[48697] == 48697 && 
b[48698] == 48698 && 
b[48699] == 48699 && 
b[48700] == 48700 && 
b[48701] == 48701 && 
b[48702] == 48702 && 
b[48703] == 48703 && 
b[48704] == 48704 && 
b[48705] == 48705 && 
b[48706] == 48706 && 
b[48707] == 48707 && 
b[48708] == 48708 && 
b[48709] == 48709 && 
b[48710] == 48710 && 
b[48711] == 48711 && 
b[48712] == 48712 && 
b[48713] == 48713 && 
b[48714] == 48714 && 
b[48715] == 48715 && 
b[48716] == 48716 && 
b[48717] == 48717 && 
b[48718] == 48718 && 
b[48719] == 48719 && 
b[48720] == 48720 && 
b[48721] == 48721 && 
b[48722] == 48722 && 
b[48723] == 48723 && 
b[48724] == 48724 && 
b[48725] == 48725 && 
b[48726] == 48726 && 
b[48727] == 48727 && 
b[48728] == 48728 && 
b[48729] == 48729 && 
b[48730] == 48730 && 
b[48731] == 48731 && 
b[48732] == 48732 && 
b[48733] == 48733 && 
b[48734] == 48734 && 
b[48735] == 48735 && 
b[48736] == 48736 && 
b[48737] == 48737 && 
b[48738] == 48738 && 
b[48739] == 48739 && 
b[48740] == 48740 && 
b[48741] == 48741 && 
b[48742] == 48742 && 
b[48743] == 48743 && 
b[48744] == 48744 && 
b[48745] == 48745 && 
b[48746] == 48746 && 
b[48747] == 48747 && 
b[48748] == 48748 && 
b[48749] == 48749 && 
b[48750] == 48750 && 
b[48751] == 48751 && 
b[48752] == 48752 && 
b[48753] == 48753 && 
b[48754] == 48754 && 
b[48755] == 48755 && 
b[48756] == 48756 && 
b[48757] == 48757 && 
b[48758] == 48758 && 
b[48759] == 48759 && 
b[48760] == 48760 && 
b[48761] == 48761 && 
b[48762] == 48762 && 
b[48763] == 48763 && 
b[48764] == 48764 && 
b[48765] == 48765 && 
b[48766] == 48766 && 
b[48767] == 48767 && 
b[48768] == 48768 && 
b[48769] == 48769 && 
b[48770] == 48770 && 
b[48771] == 48771 && 
b[48772] == 48772 && 
b[48773] == 48773 && 
b[48774] == 48774 && 
b[48775] == 48775 && 
b[48776] == 48776 && 
b[48777] == 48777 && 
b[48778] == 48778 && 
b[48779] == 48779 && 
b[48780] == 48780 && 
b[48781] == 48781 && 
b[48782] == 48782 && 
b[48783] == 48783 && 
b[48784] == 48784 && 
b[48785] == 48785 && 
b[48786] == 48786 && 
b[48787] == 48787 && 
b[48788] == 48788 && 
b[48789] == 48789 && 
b[48790] == 48790 && 
b[48791] == 48791 && 
b[48792] == 48792 && 
b[48793] == 48793 && 
b[48794] == 48794 && 
b[48795] == 48795 && 
b[48796] == 48796 && 
b[48797] == 48797 && 
b[48798] == 48798 && 
b[48799] == 48799 && 
b[48800] == 48800 && 
b[48801] == 48801 && 
b[48802] == 48802 && 
b[48803] == 48803 && 
b[48804] == 48804 && 
b[48805] == 48805 && 
b[48806] == 48806 && 
b[48807] == 48807 && 
b[48808] == 48808 && 
b[48809] == 48809 && 
b[48810] == 48810 && 
b[48811] == 48811 && 
b[48812] == 48812 && 
b[48813] == 48813 && 
b[48814] == 48814 && 
b[48815] == 48815 && 
b[48816] == 48816 && 
b[48817] == 48817 && 
b[48818] == 48818 && 
b[48819] == 48819 && 
b[48820] == 48820 && 
b[48821] == 48821 && 
b[48822] == 48822 && 
b[48823] == 48823 && 
b[48824] == 48824 && 
b[48825] == 48825 && 
b[48826] == 48826 && 
b[48827] == 48827 && 
b[48828] == 48828 && 
b[48829] == 48829 && 
b[48830] == 48830 && 
b[48831] == 48831 && 
b[48832] == 48832 && 
b[48833] == 48833 && 
b[48834] == 48834 && 
b[48835] == 48835 && 
b[48836] == 48836 && 
b[48837] == 48837 && 
b[48838] == 48838 && 
b[48839] == 48839 && 
b[48840] == 48840 && 
b[48841] == 48841 && 
b[48842] == 48842 && 
b[48843] == 48843 && 
b[48844] == 48844 && 
b[48845] == 48845 && 
b[48846] == 48846 && 
b[48847] == 48847 && 
b[48848] == 48848 && 
b[48849] == 48849 && 
b[48850] == 48850 && 
b[48851] == 48851 && 
b[48852] == 48852 && 
b[48853] == 48853 && 
b[48854] == 48854 && 
b[48855] == 48855 && 
b[48856] == 48856 && 
b[48857] == 48857 && 
b[48858] == 48858 && 
b[48859] == 48859 && 
b[48860] == 48860 && 
b[48861] == 48861 && 
b[48862] == 48862 && 
b[48863] == 48863 && 
b[48864] == 48864 && 
b[48865] == 48865 && 
b[48866] == 48866 && 
b[48867] == 48867 && 
b[48868] == 48868 && 
b[48869] == 48869 && 
b[48870] == 48870 && 
b[48871] == 48871 && 
b[48872] == 48872 && 
b[48873] == 48873 && 
b[48874] == 48874 && 
b[48875] == 48875 && 
b[48876] == 48876 && 
b[48877] == 48877 && 
b[48878] == 48878 && 
b[48879] == 48879 && 
b[48880] == 48880 && 
b[48881] == 48881 && 
b[48882] == 48882 && 
b[48883] == 48883 && 
b[48884] == 48884 && 
b[48885] == 48885 && 
b[48886] == 48886 && 
b[48887] == 48887 && 
b[48888] == 48888 && 
b[48889] == 48889 && 
b[48890] == 48890 && 
b[48891] == 48891 && 
b[48892] == 48892 && 
b[48893] == 48893 && 
b[48894] == 48894 && 
b[48895] == 48895 && 
b[48896] == 48896 && 
b[48897] == 48897 && 
b[48898] == 48898 && 
b[48899] == 48899 && 
b[48900] == 48900 && 
b[48901] == 48901 && 
b[48902] == 48902 && 
b[48903] == 48903 && 
b[48904] == 48904 && 
b[48905] == 48905 && 
b[48906] == 48906 && 
b[48907] == 48907 && 
b[48908] == 48908 && 
b[48909] == 48909 && 
b[48910] == 48910 && 
b[48911] == 48911 && 
b[48912] == 48912 && 
b[48913] == 48913 && 
b[48914] == 48914 && 
b[48915] == 48915 && 
b[48916] == 48916 && 
b[48917] == 48917 && 
b[48918] == 48918 && 
b[48919] == 48919 && 
b[48920] == 48920 && 
b[48921] == 48921 && 
b[48922] == 48922 && 
b[48923] == 48923 && 
b[48924] == 48924 && 
b[48925] == 48925 && 
b[48926] == 48926 && 
b[48927] == 48927 && 
b[48928] == 48928 && 
b[48929] == 48929 && 
b[48930] == 48930 && 
b[48931] == 48931 && 
b[48932] == 48932 && 
b[48933] == 48933 && 
b[48934] == 48934 && 
b[48935] == 48935 && 
b[48936] == 48936 && 
b[48937] == 48937 && 
b[48938] == 48938 && 
b[48939] == 48939 && 
b[48940] == 48940 && 
b[48941] == 48941 && 
b[48942] == 48942 && 
b[48943] == 48943 && 
b[48944] == 48944 && 
b[48945] == 48945 && 
b[48946] == 48946 && 
b[48947] == 48947 && 
b[48948] == 48948 && 
b[48949] == 48949 && 
b[48950] == 48950 && 
b[48951] == 48951 && 
b[48952] == 48952 && 
b[48953] == 48953 && 
b[48954] == 48954 && 
b[48955] == 48955 && 
b[48956] == 48956 && 
b[48957] == 48957 && 
b[48958] == 48958 && 
b[48959] == 48959 && 
b[48960] == 48960 && 
b[48961] == 48961 && 
b[48962] == 48962 && 
b[48963] == 48963 && 
b[48964] == 48964 && 
b[48965] == 48965 && 
b[48966] == 48966 && 
b[48967] == 48967 && 
b[48968] == 48968 && 
b[48969] == 48969 && 
b[48970] == 48970 && 
b[48971] == 48971 && 
b[48972] == 48972 && 
b[48973] == 48973 && 
b[48974] == 48974 && 
b[48975] == 48975 && 
b[48976] == 48976 && 
b[48977] == 48977 && 
b[48978] == 48978 && 
b[48979] == 48979 && 
b[48980] == 48980 && 
b[48981] == 48981 && 
b[48982] == 48982 && 
b[48983] == 48983 && 
b[48984] == 48984 && 
b[48985] == 48985 && 
b[48986] == 48986 && 
b[48987] == 48987 && 
b[48988] == 48988 && 
b[48989] == 48989 && 
b[48990] == 48990 && 
b[48991] == 48991 && 
b[48992] == 48992 && 
b[48993] == 48993 && 
b[48994] == 48994 && 
b[48995] == 48995 && 
b[48996] == 48996 && 
b[48997] == 48997 && 
b[48998] == 48998 && 
b[48999] == 48999 && 
b[49000] == 49000 && 
b[49001] == 49001 && 
b[49002] == 49002 && 
b[49003] == 49003 && 
b[49004] == 49004 && 
b[49005] == 49005 && 
b[49006] == 49006 && 
b[49007] == 49007 && 
b[49008] == 49008 && 
b[49009] == 49009 && 
b[49010] == 49010 && 
b[49011] == 49011 && 
b[49012] == 49012 && 
b[49013] == 49013 && 
b[49014] == 49014 && 
b[49015] == 49015 && 
b[49016] == 49016 && 
b[49017] == 49017 && 
b[49018] == 49018 && 
b[49019] == 49019 && 
b[49020] == 49020 && 
b[49021] == 49021 && 
b[49022] == 49022 && 
b[49023] == 49023 && 
b[49024] == 49024 && 
b[49025] == 49025 && 
b[49026] == 49026 && 
b[49027] == 49027 && 
b[49028] == 49028 && 
b[49029] == 49029 && 
b[49030] == 49030 && 
b[49031] == 49031 && 
b[49032] == 49032 && 
b[49033] == 49033 && 
b[49034] == 49034 && 
b[49035] == 49035 && 
b[49036] == 49036 && 
b[49037] == 49037 && 
b[49038] == 49038 && 
b[49039] == 49039 && 
b[49040] == 49040 && 
b[49041] == 49041 && 
b[49042] == 49042 && 
b[49043] == 49043 && 
b[49044] == 49044 && 
b[49045] == 49045 && 
b[49046] == 49046 && 
b[49047] == 49047 && 
b[49048] == 49048 && 
b[49049] == 49049 && 
b[49050] == 49050 && 
b[49051] == 49051 && 
b[49052] == 49052 && 
b[49053] == 49053 && 
b[49054] == 49054 && 
b[49055] == 49055 && 
b[49056] == 49056 && 
b[49057] == 49057 && 
b[49058] == 49058 && 
b[49059] == 49059 && 
b[49060] == 49060 && 
b[49061] == 49061 && 
b[49062] == 49062 && 
b[49063] == 49063 && 
b[49064] == 49064 && 
b[49065] == 49065 && 
b[49066] == 49066 && 
b[49067] == 49067 && 
b[49068] == 49068 && 
b[49069] == 49069 && 
b[49070] == 49070 && 
b[49071] == 49071 && 
b[49072] == 49072 && 
b[49073] == 49073 && 
b[49074] == 49074 && 
b[49075] == 49075 && 
b[49076] == 49076 && 
b[49077] == 49077 && 
b[49078] == 49078 && 
b[49079] == 49079 && 
b[49080] == 49080 && 
b[49081] == 49081 && 
b[49082] == 49082 && 
b[49083] == 49083 && 
b[49084] == 49084 && 
b[49085] == 49085 && 
b[49086] == 49086 && 
b[49087] == 49087 && 
b[49088] == 49088 && 
b[49089] == 49089 && 
b[49090] == 49090 && 
b[49091] == 49091 && 
b[49092] == 49092 && 
b[49093] == 49093 && 
b[49094] == 49094 && 
b[49095] == 49095 && 
b[49096] == 49096 && 
b[49097] == 49097 && 
b[49098] == 49098 && 
b[49099] == 49099 && 
b[49100] == 49100 && 
b[49101] == 49101 && 
b[49102] == 49102 && 
b[49103] == 49103 && 
b[49104] == 49104 && 
b[49105] == 49105 && 
b[49106] == 49106 && 
b[49107] == 49107 && 
b[49108] == 49108 && 
b[49109] == 49109 && 
b[49110] == 49110 && 
b[49111] == 49111 && 
b[49112] == 49112 && 
b[49113] == 49113 && 
b[49114] == 49114 && 
b[49115] == 49115 && 
b[49116] == 49116 && 
b[49117] == 49117 && 
b[49118] == 49118 && 
b[49119] == 49119 && 
b[49120] == 49120 && 
b[49121] == 49121 && 
b[49122] == 49122 && 
b[49123] == 49123 && 
b[49124] == 49124 && 
b[49125] == 49125 && 
b[49126] == 49126 && 
b[49127] == 49127 && 
b[49128] == 49128 && 
b[49129] == 49129 && 
b[49130] == 49130 && 
b[49131] == 49131 && 
b[49132] == 49132 && 
b[49133] == 49133 && 
b[49134] == 49134 && 
b[49135] == 49135 && 
b[49136] == 49136 && 
b[49137] == 49137 && 
b[49138] == 49138 && 
b[49139] == 49139 && 
b[49140] == 49140 && 
b[49141] == 49141 && 
b[49142] == 49142 && 
b[49143] == 49143 && 
b[49144] == 49144 && 
b[49145] == 49145 && 
b[49146] == 49146 && 
b[49147] == 49147 && 
b[49148] == 49148 && 
b[49149] == 49149 && 
b[49150] == 49150 && 
b[49151] == 49151 && 
b[49152] == 49152 && 
b[49153] == 49153 && 
b[49154] == 49154 && 
b[49155] == 49155 && 
b[49156] == 49156 && 
b[49157] == 49157 && 
b[49158] == 49158 && 
b[49159] == 49159 && 
b[49160] == 49160 && 
b[49161] == 49161 && 
b[49162] == 49162 && 
b[49163] == 49163 && 
b[49164] == 49164 && 
b[49165] == 49165 && 
b[49166] == 49166 && 
b[49167] == 49167 && 
b[49168] == 49168 && 
b[49169] == 49169 && 
b[49170] == 49170 && 
b[49171] == 49171 && 
b[49172] == 49172 && 
b[49173] == 49173 && 
b[49174] == 49174 && 
b[49175] == 49175 && 
b[49176] == 49176 && 
b[49177] == 49177 && 
b[49178] == 49178 && 
b[49179] == 49179 && 
b[49180] == 49180 && 
b[49181] == 49181 && 
b[49182] == 49182 && 
b[49183] == 49183 && 
b[49184] == 49184 && 
b[49185] == 49185 && 
b[49186] == 49186 && 
b[49187] == 49187 && 
b[49188] == 49188 && 
b[49189] == 49189 && 
b[49190] == 49190 && 
b[49191] == 49191 && 
b[49192] == 49192 && 
b[49193] == 49193 && 
b[49194] == 49194 && 
b[49195] == 49195 && 
b[49196] == 49196 && 
b[49197] == 49197 && 
b[49198] == 49198 && 
b[49199] == 49199 && 
b[49200] == 49200 && 
b[49201] == 49201 && 
b[49202] == 49202 && 
b[49203] == 49203 && 
b[49204] == 49204 && 
b[49205] == 49205 && 
b[49206] == 49206 && 
b[49207] == 49207 && 
b[49208] == 49208 && 
b[49209] == 49209 && 
b[49210] == 49210 && 
b[49211] == 49211 && 
b[49212] == 49212 && 
b[49213] == 49213 && 
b[49214] == 49214 && 
b[49215] == 49215 && 
b[49216] == 49216 && 
b[49217] == 49217 && 
b[49218] == 49218 && 
b[49219] == 49219 && 
b[49220] == 49220 && 
b[49221] == 49221 && 
b[49222] == 49222 && 
b[49223] == 49223 && 
b[49224] == 49224 && 
b[49225] == 49225 && 
b[49226] == 49226 && 
b[49227] == 49227 && 
b[49228] == 49228 && 
b[49229] == 49229 && 
b[49230] == 49230 && 
b[49231] == 49231 && 
b[49232] == 49232 && 
b[49233] == 49233 && 
b[49234] == 49234 && 
b[49235] == 49235 && 
b[49236] == 49236 && 
b[49237] == 49237 && 
b[49238] == 49238 && 
b[49239] == 49239 && 
b[49240] == 49240 && 
b[49241] == 49241 && 
b[49242] == 49242 && 
b[49243] == 49243 && 
b[49244] == 49244 && 
b[49245] == 49245 && 
b[49246] == 49246 && 
b[49247] == 49247 && 
b[49248] == 49248 && 
b[49249] == 49249 && 
b[49250] == 49250 && 
b[49251] == 49251 && 
b[49252] == 49252 && 
b[49253] == 49253 && 
b[49254] == 49254 && 
b[49255] == 49255 && 
b[49256] == 49256 && 
b[49257] == 49257 && 
b[49258] == 49258 && 
b[49259] == 49259 && 
b[49260] == 49260 && 
b[49261] == 49261 && 
b[49262] == 49262 && 
b[49263] == 49263 && 
b[49264] == 49264 && 
b[49265] == 49265 && 
b[49266] == 49266 && 
b[49267] == 49267 && 
b[49268] == 49268 && 
b[49269] == 49269 && 
b[49270] == 49270 && 
b[49271] == 49271 && 
b[49272] == 49272 && 
b[49273] == 49273 && 
b[49274] == 49274 && 
b[49275] == 49275 && 
b[49276] == 49276 && 
b[49277] == 49277 && 
b[49278] == 49278 && 
b[49279] == 49279 && 
b[49280] == 49280 && 
b[49281] == 49281 && 
b[49282] == 49282 && 
b[49283] == 49283 && 
b[49284] == 49284 && 
b[49285] == 49285 && 
b[49286] == 49286 && 
b[49287] == 49287 && 
b[49288] == 49288 && 
b[49289] == 49289 && 
b[49290] == 49290 && 
b[49291] == 49291 && 
b[49292] == 49292 && 
b[49293] == 49293 && 
b[49294] == 49294 && 
b[49295] == 49295 && 
b[49296] == 49296 && 
b[49297] == 49297 && 
b[49298] == 49298 && 
b[49299] == 49299 && 
b[49300] == 49300 && 
b[49301] == 49301 && 
b[49302] == 49302 && 
b[49303] == 49303 && 
b[49304] == 49304 && 
b[49305] == 49305 && 
b[49306] == 49306 && 
b[49307] == 49307 && 
b[49308] == 49308 && 
b[49309] == 49309 && 
b[49310] == 49310 && 
b[49311] == 49311 && 
b[49312] == 49312 && 
b[49313] == 49313 && 
b[49314] == 49314 && 
b[49315] == 49315 && 
b[49316] == 49316 && 
b[49317] == 49317 && 
b[49318] == 49318 && 
b[49319] == 49319 && 
b[49320] == 49320 && 
b[49321] == 49321 && 
b[49322] == 49322 && 
b[49323] == 49323 && 
b[49324] == 49324 && 
b[49325] == 49325 && 
b[49326] == 49326 && 
b[49327] == 49327 && 
b[49328] == 49328 && 
b[49329] == 49329 && 
b[49330] == 49330 && 
b[49331] == 49331 && 
b[49332] == 49332 && 
b[49333] == 49333 && 
b[49334] == 49334 && 
b[49335] == 49335 && 
b[49336] == 49336 && 
b[49337] == 49337 && 
b[49338] == 49338 && 
b[49339] == 49339 && 
b[49340] == 49340 && 
b[49341] == 49341 && 
b[49342] == 49342 && 
b[49343] == 49343 && 
b[49344] == 49344 && 
b[49345] == 49345 && 
b[49346] == 49346 && 
b[49347] == 49347 && 
b[49348] == 49348 && 
b[49349] == 49349 && 
b[49350] == 49350 && 
b[49351] == 49351 && 
b[49352] == 49352 && 
b[49353] == 49353 && 
b[49354] == 49354 && 
b[49355] == 49355 && 
b[49356] == 49356 && 
b[49357] == 49357 && 
b[49358] == 49358 && 
b[49359] == 49359 && 
b[49360] == 49360 && 
b[49361] == 49361 && 
b[49362] == 49362 && 
b[49363] == 49363 && 
b[49364] == 49364 && 
b[49365] == 49365 && 
b[49366] == 49366 && 
b[49367] == 49367 && 
b[49368] == 49368 && 
b[49369] == 49369 && 
b[49370] == 49370 && 
b[49371] == 49371 && 
b[49372] == 49372 && 
b[49373] == 49373 && 
b[49374] == 49374 && 
b[49375] == 49375 && 
b[49376] == 49376 && 
b[49377] == 49377 && 
b[49378] == 49378 && 
b[49379] == 49379 && 
b[49380] == 49380 && 
b[49381] == 49381 && 
b[49382] == 49382 && 
b[49383] == 49383 && 
b[49384] == 49384 && 
b[49385] == 49385 && 
b[49386] == 49386 && 
b[49387] == 49387 && 
b[49388] == 49388 && 
b[49389] == 49389 && 
b[49390] == 49390 && 
b[49391] == 49391 && 
b[49392] == 49392 && 
b[49393] == 49393 && 
b[49394] == 49394 && 
b[49395] == 49395 && 
b[49396] == 49396 && 
b[49397] == 49397 && 
b[49398] == 49398 && 
b[49399] == 49399 && 
b[49400] == 49400 && 
b[49401] == 49401 && 
b[49402] == 49402 && 
b[49403] == 49403 && 
b[49404] == 49404 && 
b[49405] == 49405 && 
b[49406] == 49406 && 
b[49407] == 49407 && 
b[49408] == 49408 && 
b[49409] == 49409 && 
b[49410] == 49410 && 
b[49411] == 49411 && 
b[49412] == 49412 && 
b[49413] == 49413 && 
b[49414] == 49414 && 
b[49415] == 49415 && 
b[49416] == 49416 && 
b[49417] == 49417 && 
b[49418] == 49418 && 
b[49419] == 49419 && 
b[49420] == 49420 && 
b[49421] == 49421 && 
b[49422] == 49422 && 
b[49423] == 49423 && 
b[49424] == 49424 && 
b[49425] == 49425 && 
b[49426] == 49426 && 
b[49427] == 49427 && 
b[49428] == 49428 && 
b[49429] == 49429 && 
b[49430] == 49430 && 
b[49431] == 49431 && 
b[49432] == 49432 && 
b[49433] == 49433 && 
b[49434] == 49434 && 
b[49435] == 49435 && 
b[49436] == 49436 && 
b[49437] == 49437 && 
b[49438] == 49438 && 
b[49439] == 49439 && 
b[49440] == 49440 && 
b[49441] == 49441 && 
b[49442] == 49442 && 
b[49443] == 49443 && 
b[49444] == 49444 && 
b[49445] == 49445 && 
b[49446] == 49446 && 
b[49447] == 49447 && 
b[49448] == 49448 && 
b[49449] == 49449 && 
b[49450] == 49450 && 
b[49451] == 49451 && 
b[49452] == 49452 && 
b[49453] == 49453 && 
b[49454] == 49454 && 
b[49455] == 49455 && 
b[49456] == 49456 && 
b[49457] == 49457 && 
b[49458] == 49458 && 
b[49459] == 49459 && 
b[49460] == 49460 && 
b[49461] == 49461 && 
b[49462] == 49462 && 
b[49463] == 49463 && 
b[49464] == 49464 && 
b[49465] == 49465 && 
b[49466] == 49466 && 
b[49467] == 49467 && 
b[49468] == 49468 && 
b[49469] == 49469 && 
b[49470] == 49470 && 
b[49471] == 49471 && 
b[49472] == 49472 && 
b[49473] == 49473 && 
b[49474] == 49474 && 
b[49475] == 49475 && 
b[49476] == 49476 && 
b[49477] == 49477 && 
b[49478] == 49478 && 
b[49479] == 49479 && 
b[49480] == 49480 && 
b[49481] == 49481 && 
b[49482] == 49482 && 
b[49483] == 49483 && 
b[49484] == 49484 && 
b[49485] == 49485 && 
b[49486] == 49486 && 
b[49487] == 49487 && 
b[49488] == 49488 && 
b[49489] == 49489 && 
b[49490] == 49490 && 
b[49491] == 49491 && 
b[49492] == 49492 && 
b[49493] == 49493 && 
b[49494] == 49494 && 
b[49495] == 49495 && 
b[49496] == 49496 && 
b[49497] == 49497 && 
b[49498] == 49498 && 
b[49499] == 49499 && 
b[49500] == 49500 && 
b[49501] == 49501 && 
b[49502] == 49502 && 
b[49503] == 49503 && 
b[49504] == 49504 && 
b[49505] == 49505 && 
b[49506] == 49506 && 
b[49507] == 49507 && 
b[49508] == 49508 && 
b[49509] == 49509 && 
b[49510] == 49510 && 
b[49511] == 49511 && 
b[49512] == 49512 && 
b[49513] == 49513 && 
b[49514] == 49514 && 
b[49515] == 49515 && 
b[49516] == 49516 && 
b[49517] == 49517 && 
b[49518] == 49518 && 
b[49519] == 49519 && 
b[49520] == 49520 && 
b[49521] == 49521 && 
b[49522] == 49522 && 
b[49523] == 49523 && 
b[49524] == 49524 && 
b[49525] == 49525 && 
b[49526] == 49526 && 
b[49527] == 49527 && 
b[49528] == 49528 && 
b[49529] == 49529 && 
b[49530] == 49530 && 
b[49531] == 49531 && 
b[49532] == 49532 && 
b[49533] == 49533 && 
b[49534] == 49534 && 
b[49535] == 49535 && 
b[49536] == 49536 && 
b[49537] == 49537 && 
b[49538] == 49538 && 
b[49539] == 49539 && 
b[49540] == 49540 && 
b[49541] == 49541 && 
b[49542] == 49542 && 
b[49543] == 49543 && 
b[49544] == 49544 && 
b[49545] == 49545 && 
b[49546] == 49546 && 
b[49547] == 49547 && 
b[49548] == 49548 && 
b[49549] == 49549 && 
b[49550] == 49550 && 
b[49551] == 49551 && 
b[49552] == 49552 && 
b[49553] == 49553 && 
b[49554] == 49554 && 
b[49555] == 49555 && 
b[49556] == 49556 && 
b[49557] == 49557 && 
b[49558] == 49558 && 
b[49559] == 49559 && 
b[49560] == 49560 && 
b[49561] == 49561 && 
b[49562] == 49562 && 
b[49563] == 49563 && 
b[49564] == 49564 && 
b[49565] == 49565 && 
b[49566] == 49566 && 
b[49567] == 49567 && 
b[49568] == 49568 && 
b[49569] == 49569 && 
b[49570] == 49570 && 
b[49571] == 49571 && 
b[49572] == 49572 && 
b[49573] == 49573 && 
b[49574] == 49574 && 
b[49575] == 49575 && 
b[49576] == 49576 && 
b[49577] == 49577 && 
b[49578] == 49578 && 
b[49579] == 49579 && 
b[49580] == 49580 && 
b[49581] == 49581 && 
b[49582] == 49582 && 
b[49583] == 49583 && 
b[49584] == 49584 && 
b[49585] == 49585 && 
b[49586] == 49586 && 
b[49587] == 49587 && 
b[49588] == 49588 && 
b[49589] == 49589 && 
b[49590] == 49590 && 
b[49591] == 49591 && 
b[49592] == 49592 && 
b[49593] == 49593 && 
b[49594] == 49594 && 
b[49595] == 49595 && 
b[49596] == 49596 && 
b[49597] == 49597 && 
b[49598] == 49598 && 
b[49599] == 49599 && 
b[49600] == 49600 && 
b[49601] == 49601 && 
b[49602] == 49602 && 
b[49603] == 49603 && 
b[49604] == 49604 && 
b[49605] == 49605 && 
b[49606] == 49606 && 
b[49607] == 49607 && 
b[49608] == 49608 && 
b[49609] == 49609 && 
b[49610] == 49610 && 
b[49611] == 49611 && 
b[49612] == 49612 && 
b[49613] == 49613 && 
b[49614] == 49614 && 
b[49615] == 49615 && 
b[49616] == 49616 && 
b[49617] == 49617 && 
b[49618] == 49618 && 
b[49619] == 49619 && 
b[49620] == 49620 && 
b[49621] == 49621 && 
b[49622] == 49622 && 
b[49623] == 49623 && 
b[49624] == 49624 && 
b[49625] == 49625 && 
b[49626] == 49626 && 
b[49627] == 49627 && 
b[49628] == 49628 && 
b[49629] == 49629 && 
b[49630] == 49630 && 
b[49631] == 49631 && 
b[49632] == 49632 && 
b[49633] == 49633 && 
b[49634] == 49634 && 
b[49635] == 49635 && 
b[49636] == 49636 && 
b[49637] == 49637 && 
b[49638] == 49638 && 
b[49639] == 49639 && 
b[49640] == 49640 && 
b[49641] == 49641 && 
b[49642] == 49642 && 
b[49643] == 49643 && 
b[49644] == 49644 && 
b[49645] == 49645 && 
b[49646] == 49646 && 
b[49647] == 49647 && 
b[49648] == 49648 && 
b[49649] == 49649 && 
b[49650] == 49650 && 
b[49651] == 49651 && 
b[49652] == 49652 && 
b[49653] == 49653 && 
b[49654] == 49654 && 
b[49655] == 49655 && 
b[49656] == 49656 && 
b[49657] == 49657 && 
b[49658] == 49658 && 
b[49659] == 49659 && 
b[49660] == 49660 && 
b[49661] == 49661 && 
b[49662] == 49662 && 
b[49663] == 49663 && 
b[49664] == 49664 && 
b[49665] == 49665 && 
b[49666] == 49666 && 
b[49667] == 49667 && 
b[49668] == 49668 && 
b[49669] == 49669 && 
b[49670] == 49670 && 
b[49671] == 49671 && 
b[49672] == 49672 && 
b[49673] == 49673 && 
b[49674] == 49674 && 
b[49675] == 49675 && 
b[49676] == 49676 && 
b[49677] == 49677 && 
b[49678] == 49678 && 
b[49679] == 49679 && 
b[49680] == 49680 && 
b[49681] == 49681 && 
b[49682] == 49682 && 
b[49683] == 49683 && 
b[49684] == 49684 && 
b[49685] == 49685 && 
b[49686] == 49686 && 
b[49687] == 49687 && 
b[49688] == 49688 && 
b[49689] == 49689 && 
b[49690] == 49690 && 
b[49691] == 49691 && 
b[49692] == 49692 && 
b[49693] == 49693 && 
b[49694] == 49694 && 
b[49695] == 49695 && 
b[49696] == 49696 && 
b[49697] == 49697 && 
b[49698] == 49698 && 
b[49699] == 49699 && 
b[49700] == 49700 && 
b[49701] == 49701 && 
b[49702] == 49702 && 
b[49703] == 49703 && 
b[49704] == 49704 && 
b[49705] == 49705 && 
b[49706] == 49706 && 
b[49707] == 49707 && 
b[49708] == 49708 && 
b[49709] == 49709 && 
b[49710] == 49710 && 
b[49711] == 49711 && 
b[49712] == 49712 && 
b[49713] == 49713 && 
b[49714] == 49714 && 
b[49715] == 49715 && 
b[49716] == 49716 && 
b[49717] == 49717 && 
b[49718] == 49718 && 
b[49719] == 49719 && 
b[49720] == 49720 && 
b[49721] == 49721 && 
b[49722] == 49722 && 
b[49723] == 49723 && 
b[49724] == 49724 && 
b[49725] == 49725 && 
b[49726] == 49726 && 
b[49727] == 49727 && 
b[49728] == 49728 && 
b[49729] == 49729 && 
b[49730] == 49730 && 
b[49731] == 49731 && 
b[49732] == 49732 && 
b[49733] == 49733 && 
b[49734] == 49734 && 
b[49735] == 49735 && 
b[49736] == 49736 && 
b[49737] == 49737 && 
b[49738] == 49738 && 
b[49739] == 49739 && 
b[49740] == 49740 && 
b[49741] == 49741 && 
b[49742] == 49742 && 
b[49743] == 49743 && 
b[49744] == 49744 && 
b[49745] == 49745 && 
b[49746] == 49746 && 
b[49747] == 49747 && 
b[49748] == 49748 && 
b[49749] == 49749 && 
b[49750] == 49750 && 
b[49751] == 49751 && 
b[49752] == 49752 && 
b[49753] == 49753 && 
b[49754] == 49754 && 
b[49755] == 49755 && 
b[49756] == 49756 && 
b[49757] == 49757 && 
b[49758] == 49758 && 
b[49759] == 49759 && 
b[49760] == 49760 && 
b[49761] == 49761 && 
b[49762] == 49762 && 
b[49763] == 49763 && 
b[49764] == 49764 && 
b[49765] == 49765 && 
b[49766] == 49766 && 
b[49767] == 49767 && 
b[49768] == 49768 && 
b[49769] == 49769 && 
b[49770] == 49770 && 
b[49771] == 49771 && 
b[49772] == 49772 && 
b[49773] == 49773 && 
b[49774] == 49774 && 
b[49775] == 49775 && 
b[49776] == 49776 && 
b[49777] == 49777 && 
b[49778] == 49778 && 
b[49779] == 49779 && 
b[49780] == 49780 && 
b[49781] == 49781 && 
b[49782] == 49782 && 
b[49783] == 49783 && 
b[49784] == 49784 && 
b[49785] == 49785 && 
b[49786] == 49786 && 
b[49787] == 49787 && 
b[49788] == 49788 && 
b[49789] == 49789 && 
b[49790] == 49790 && 
b[49791] == 49791 && 
b[49792] == 49792 && 
b[49793] == 49793 && 
b[49794] == 49794 && 
b[49795] == 49795 && 
b[49796] == 49796 && 
b[49797] == 49797 && 
b[49798] == 49798 && 
b[49799] == 49799 && 
b[49800] == 49800 && 
b[49801] == 49801 && 
b[49802] == 49802 && 
b[49803] == 49803 && 
b[49804] == 49804 && 
b[49805] == 49805 && 
b[49806] == 49806 && 
b[49807] == 49807 && 
b[49808] == 49808 && 
b[49809] == 49809 && 
b[49810] == 49810 && 
b[49811] == 49811 && 
b[49812] == 49812 && 
b[49813] == 49813 && 
b[49814] == 49814 && 
b[49815] == 49815 && 
b[49816] == 49816 && 
b[49817] == 49817 && 
b[49818] == 49818 && 
b[49819] == 49819 && 
b[49820] == 49820 && 
b[49821] == 49821 && 
b[49822] == 49822 && 
b[49823] == 49823 && 
b[49824] == 49824 && 
b[49825] == 49825 && 
b[49826] == 49826 && 
b[49827] == 49827 && 
b[49828] == 49828 && 
b[49829] == 49829 && 
b[49830] == 49830 && 
b[49831] == 49831 && 
b[49832] == 49832 && 
b[49833] == 49833 && 
b[49834] == 49834 && 
b[49835] == 49835 && 
b[49836] == 49836 && 
b[49837] == 49837 && 
b[49838] == 49838 && 
b[49839] == 49839 && 
b[49840] == 49840 && 
b[49841] == 49841 && 
b[49842] == 49842 && 
b[49843] == 49843 && 
b[49844] == 49844 && 
b[49845] == 49845 && 
b[49846] == 49846 && 
b[49847] == 49847 && 
b[49848] == 49848 && 
b[49849] == 49849 && 
b[49850] == 49850 && 
b[49851] == 49851 && 
b[49852] == 49852 && 
b[49853] == 49853 && 
b[49854] == 49854 && 
b[49855] == 49855 && 
b[49856] == 49856 && 
b[49857] == 49857 && 
b[49858] == 49858 && 
b[49859] == 49859 && 
b[49860] == 49860 && 
b[49861] == 49861 && 
b[49862] == 49862 && 
b[49863] == 49863 && 
b[49864] == 49864 && 
b[49865] == 49865 && 
b[49866] == 49866 && 
b[49867] == 49867 && 
b[49868] == 49868 && 
b[49869] == 49869 && 
b[49870] == 49870 && 
b[49871] == 49871 && 
b[49872] == 49872 && 
b[49873] == 49873 && 
b[49874] == 49874 && 
b[49875] == 49875 && 
b[49876] == 49876 && 
b[49877] == 49877 && 
b[49878] == 49878 && 
b[49879] == 49879 && 
b[49880] == 49880 && 
b[49881] == 49881 && 
b[49882] == 49882 && 
b[49883] == 49883 && 
b[49884] == 49884 && 
b[49885] == 49885 && 
b[49886] == 49886 && 
b[49887] == 49887 && 
b[49888] == 49888 && 
b[49889] == 49889 && 
b[49890] == 49890 && 
b[49891] == 49891 && 
b[49892] == 49892 && 
b[49893] == 49893 && 
b[49894] == 49894 && 
b[49895] == 49895 && 
b[49896] == 49896 && 
b[49897] == 49897 && 
b[49898] == 49898 && 
b[49899] == 49899 && 
b[49900] == 49900 && 
b[49901] == 49901 && 
b[49902] == 49902 && 
b[49903] == 49903 && 
b[49904] == 49904 && 
b[49905] == 49905 && 
b[49906] == 49906 && 
b[49907] == 49907 && 
b[49908] == 49908 && 
b[49909] == 49909 && 
b[49910] == 49910 && 
b[49911] == 49911 && 
b[49912] == 49912 && 
b[49913] == 49913 && 
b[49914] == 49914 && 
b[49915] == 49915 && 
b[49916] == 49916 && 
b[49917] == 49917 && 
b[49918] == 49918 && 
b[49919] == 49919 && 
b[49920] == 49920 && 
b[49921] == 49921 && 
b[49922] == 49922 && 
b[49923] == 49923 && 
b[49924] == 49924 && 
b[49925] == 49925 && 
b[49926] == 49926 && 
b[49927] == 49927 && 
b[49928] == 49928 && 
b[49929] == 49929 && 
b[49930] == 49930 && 
b[49931] == 49931 && 
b[49932] == 49932 && 
b[49933] == 49933 && 
b[49934] == 49934 && 
b[49935] == 49935 && 
b[49936] == 49936 && 
b[49937] == 49937 && 
b[49938] == 49938 && 
b[49939] == 49939 && 
b[49940] == 49940 && 
b[49941] == 49941 && 
b[49942] == 49942 && 
b[49943] == 49943 && 
b[49944] == 49944 && 
b[49945] == 49945 && 
b[49946] == 49946 && 
b[49947] == 49947 && 
b[49948] == 49948 && 
b[49949] == 49949 && 
b[49950] == 49950 && 
b[49951] == 49951 && 
b[49952] == 49952 && 
b[49953] == 49953 && 
b[49954] == 49954 && 
b[49955] == 49955 && 
b[49956] == 49956 && 
b[49957] == 49957 && 
b[49958] == 49958 && 
b[49959] == 49959 && 
b[49960] == 49960 && 
b[49961] == 49961 && 
b[49962] == 49962 && 
b[49963] == 49963 && 
b[49964] == 49964 && 
b[49965] == 49965 && 
b[49966] == 49966 && 
b[49967] == 49967 && 
b[49968] == 49968 && 
b[49969] == 49969 && 
b[49970] == 49970 && 
b[49971] == 49971 && 
b[49972] == 49972 && 
b[49973] == 49973 && 
b[49974] == 49974 && 
b[49975] == 49975 && 
b[49976] == 49976 && 
b[49977] == 49977 && 
b[49978] == 49978 && 
b[49979] == 49979 && 
b[49980] == 49980 && 
b[49981] == 49981 && 
b[49982] == 49982 && 
b[49983] == 49983 && 
b[49984] == 49984 && 
b[49985] == 49985 && 
b[49986] == 49986 && 
b[49987] == 49987 && 
b[49988] == 49988 && 
b[49989] == 49989 && 
b[49990] == 49990 && 
b[49991] == 49991 && 
b[49992] == 49992 && 
b[49993] == 49993 && 
b[49994] == 49994 && 
b[49995] == 49995 && 
b[49996] == 49996 && 
b[49997] == 49997 && 
b[49998] == 49998 && 
b[49999] == 49999 && 
b[50000] == 50000 && 
b[50001] == 50001 && 
b[50002] == 50002 && 
b[50003] == 50003 && 
b[50004] == 50004 && 
b[50005] == 50005 && 
b[50006] == 50006 && 
b[50007] == 50007 && 
b[50008] == 50008 && 
b[50009] == 50009 && 
b[50010] == 50010 && 
b[50011] == 50011 && 
b[50012] == 50012 && 
b[50013] == 50013 && 
b[50014] == 50014 && 
b[50015] == 50015 && 
b[50016] == 50016 && 
b[50017] == 50017 && 
b[50018] == 50018 && 
b[50019] == 50019 && 
b[50020] == 50020 && 
b[50021] == 50021 && 
b[50022] == 50022 && 
b[50023] == 50023 && 
b[50024] == 50024 && 
b[50025] == 50025 && 
b[50026] == 50026 && 
b[50027] == 50027 && 
b[50028] == 50028 && 
b[50029] == 50029 && 
b[50030] == 50030 && 
b[50031] == 50031 && 
b[50032] == 50032 && 
b[50033] == 50033 && 
b[50034] == 50034 && 
b[50035] == 50035 && 
b[50036] == 50036 && 
b[50037] == 50037 && 
b[50038] == 50038 && 
b[50039] == 50039 && 
b[50040] == 50040 && 
b[50041] == 50041 && 
b[50042] == 50042 && 
b[50043] == 50043 && 
b[50044] == 50044 && 
b[50045] == 50045 && 
b[50046] == 50046 && 
b[50047] == 50047 && 
b[50048] == 50048 && 
b[50049] == 50049 && 
b[50050] == 50050 && 
b[50051] == 50051 && 
b[50052] == 50052 && 
b[50053] == 50053 && 
b[50054] == 50054 && 
b[50055] == 50055 && 
b[50056] == 50056 && 
b[50057] == 50057 && 
b[50058] == 50058 && 
b[50059] == 50059 && 
b[50060] == 50060 && 
b[50061] == 50061 && 
b[50062] == 50062 && 
b[50063] == 50063 && 
b[50064] == 50064 && 
b[50065] == 50065 && 
b[50066] == 50066 && 
b[50067] == 50067 && 
b[50068] == 50068 && 
b[50069] == 50069 && 
b[50070] == 50070 && 
b[50071] == 50071 && 
b[50072] == 50072 && 
b[50073] == 50073 && 
b[50074] == 50074 && 
b[50075] == 50075 && 
b[50076] == 50076 && 
b[50077] == 50077 && 
b[50078] == 50078 && 
b[50079] == 50079 && 
b[50080] == 50080 && 
b[50081] == 50081 && 
b[50082] == 50082 && 
b[50083] == 50083 && 
b[50084] == 50084 && 
b[50085] == 50085 && 
b[50086] == 50086 && 
b[50087] == 50087 && 
b[50088] == 50088 && 
b[50089] == 50089 && 
b[50090] == 50090 && 
b[50091] == 50091 && 
b[50092] == 50092 && 
b[50093] == 50093 && 
b[50094] == 50094 && 
b[50095] == 50095 && 
b[50096] == 50096 && 
b[50097] == 50097 && 
b[50098] == 50098 && 
b[50099] == 50099 && 
b[50100] == 50100 && 
b[50101] == 50101 && 
b[50102] == 50102 && 
b[50103] == 50103 && 
b[50104] == 50104 && 
b[50105] == 50105 && 
b[50106] == 50106 && 
b[50107] == 50107 && 
b[50108] == 50108 && 
b[50109] == 50109 && 
b[50110] == 50110 && 
b[50111] == 50111 && 
b[50112] == 50112 && 
b[50113] == 50113 && 
b[50114] == 50114 && 
b[50115] == 50115 && 
b[50116] == 50116 && 
b[50117] == 50117 && 
b[50118] == 50118 && 
b[50119] == 50119 && 
b[50120] == 50120 && 
b[50121] == 50121 && 
b[50122] == 50122 && 
b[50123] == 50123 && 
b[50124] == 50124 && 
b[50125] == 50125 && 
b[50126] == 50126 && 
b[50127] == 50127 && 
b[50128] == 50128 && 
b[50129] == 50129 && 
b[50130] == 50130 && 
b[50131] == 50131 && 
b[50132] == 50132 && 
b[50133] == 50133 && 
b[50134] == 50134 && 
b[50135] == 50135 && 
b[50136] == 50136 && 
b[50137] == 50137 && 
b[50138] == 50138 && 
b[50139] == 50139 && 
b[50140] == 50140 && 
b[50141] == 50141 && 
b[50142] == 50142 && 
b[50143] == 50143 && 
b[50144] == 50144 && 
b[50145] == 50145 && 
b[50146] == 50146 && 
b[50147] == 50147 && 
b[50148] == 50148 && 
b[50149] == 50149 && 
b[50150] == 50150 && 
b[50151] == 50151 && 
b[50152] == 50152 && 
b[50153] == 50153 && 
b[50154] == 50154 && 
b[50155] == 50155 && 
b[50156] == 50156 && 
b[50157] == 50157 && 
b[50158] == 50158 && 
b[50159] == 50159 && 
b[50160] == 50160 && 
b[50161] == 50161 && 
b[50162] == 50162 && 
b[50163] == 50163 && 
b[50164] == 50164 && 
b[50165] == 50165 && 
b[50166] == 50166 && 
b[50167] == 50167 && 
b[50168] == 50168 && 
b[50169] == 50169 && 
b[50170] == 50170 && 
b[50171] == 50171 && 
b[50172] == 50172 && 
b[50173] == 50173 && 
b[50174] == 50174 && 
b[50175] == 50175 && 
b[50176] == 50176 && 
b[50177] == 50177 && 
b[50178] == 50178 && 
b[50179] == 50179 && 
b[50180] == 50180 && 
b[50181] == 50181 && 
b[50182] == 50182 && 
b[50183] == 50183 && 
b[50184] == 50184 && 
b[50185] == 50185 && 
b[50186] == 50186 && 
b[50187] == 50187 && 
b[50188] == 50188 && 
b[50189] == 50189 && 
b[50190] == 50190 && 
b[50191] == 50191 && 
b[50192] == 50192 && 
b[50193] == 50193 && 
b[50194] == 50194 && 
b[50195] == 50195 && 
b[50196] == 50196 && 
b[50197] == 50197 && 
b[50198] == 50198 && 
b[50199] == 50199 && 
b[50200] == 50200 && 
b[50201] == 50201 && 
b[50202] == 50202 && 
b[50203] == 50203 && 
b[50204] == 50204 && 
b[50205] == 50205 && 
b[50206] == 50206 && 
b[50207] == 50207 && 
b[50208] == 50208 && 
b[50209] == 50209 && 
b[50210] == 50210 && 
b[50211] == 50211 && 
b[50212] == 50212 && 
b[50213] == 50213 && 
b[50214] == 50214 && 
b[50215] == 50215 && 
b[50216] == 50216 && 
b[50217] == 50217 && 
b[50218] == 50218 && 
b[50219] == 50219 && 
b[50220] == 50220 && 
b[50221] == 50221 && 
b[50222] == 50222 && 
b[50223] == 50223 && 
b[50224] == 50224 && 
b[50225] == 50225 && 
b[50226] == 50226 && 
b[50227] == 50227 && 
b[50228] == 50228 && 
b[50229] == 50229 && 
b[50230] == 50230 && 
b[50231] == 50231 && 
b[50232] == 50232 && 
b[50233] == 50233 && 
b[50234] == 50234 && 
b[50235] == 50235 && 
b[50236] == 50236 && 
b[50237] == 50237 && 
b[50238] == 50238 && 
b[50239] == 50239 && 
b[50240] == 50240 && 
b[50241] == 50241 && 
b[50242] == 50242 && 
b[50243] == 50243 && 
b[50244] == 50244 && 
b[50245] == 50245 && 
b[50246] == 50246 && 
b[50247] == 50247 && 
b[50248] == 50248 && 
b[50249] == 50249 && 
b[50250] == 50250 && 
b[50251] == 50251 && 
b[50252] == 50252 && 
b[50253] == 50253 && 
b[50254] == 50254 && 
b[50255] == 50255 && 
b[50256] == 50256 && 
b[50257] == 50257 && 
b[50258] == 50258 && 
b[50259] == 50259 && 
b[50260] == 50260 && 
b[50261] == 50261 && 
b[50262] == 50262 && 
b[50263] == 50263 && 
b[50264] == 50264 && 
b[50265] == 50265 && 
b[50266] == 50266 && 
b[50267] == 50267 && 
b[50268] == 50268 && 
b[50269] == 50269 && 
b[50270] == 50270 && 
b[50271] == 50271 && 
b[50272] == 50272 && 
b[50273] == 50273 && 
b[50274] == 50274 && 
b[50275] == 50275 && 
b[50276] == 50276 && 
b[50277] == 50277 && 
b[50278] == 50278 && 
b[50279] == 50279 && 
b[50280] == 50280 && 
b[50281] == 50281 && 
b[50282] == 50282 && 
b[50283] == 50283 && 
b[50284] == 50284 && 
b[50285] == 50285 && 
b[50286] == 50286 && 
b[50287] == 50287 && 
b[50288] == 50288 && 
b[50289] == 50289 && 
b[50290] == 50290 && 
b[50291] == 50291 && 
b[50292] == 50292 && 
b[50293] == 50293 && 
b[50294] == 50294 && 
b[50295] == 50295 && 
b[50296] == 50296 && 
b[50297] == 50297 && 
b[50298] == 50298 && 
b[50299] == 50299 && 
b[50300] == 50300 && 
b[50301] == 50301 && 
b[50302] == 50302 && 
b[50303] == 50303 && 
b[50304] == 50304 && 
b[50305] == 50305 && 
b[50306] == 50306 && 
b[50307] == 50307 && 
b[50308] == 50308 && 
b[50309] == 50309 && 
b[50310] == 50310 && 
b[50311] == 50311 && 
b[50312] == 50312 && 
b[50313] == 50313 && 
b[50314] == 50314 && 
b[50315] == 50315 && 
b[50316] == 50316 && 
b[50317] == 50317 && 
b[50318] == 50318 && 
b[50319] == 50319 && 
b[50320] == 50320 && 
b[50321] == 50321 && 
b[50322] == 50322 && 
b[50323] == 50323 && 
b[50324] == 50324 && 
b[50325] == 50325 && 
b[50326] == 50326 && 
b[50327] == 50327 && 
b[50328] == 50328 && 
b[50329] == 50329 && 
b[50330] == 50330 && 
b[50331] == 50331 && 
b[50332] == 50332 && 
b[50333] == 50333 && 
b[50334] == 50334 && 
b[50335] == 50335 && 
b[50336] == 50336 && 
b[50337] == 50337 && 
b[50338] == 50338 && 
b[50339] == 50339 && 
b[50340] == 50340 && 
b[50341] == 50341 && 
b[50342] == 50342 && 
b[50343] == 50343 && 
b[50344] == 50344 && 
b[50345] == 50345 && 
b[50346] == 50346 && 
b[50347] == 50347 && 
b[50348] == 50348 && 
b[50349] == 50349 && 
b[50350] == 50350 && 
b[50351] == 50351 && 
b[50352] == 50352 && 
b[50353] == 50353 && 
b[50354] == 50354 && 
b[50355] == 50355 && 
b[50356] == 50356 && 
b[50357] == 50357 && 
b[50358] == 50358 && 
b[50359] == 50359 && 
b[50360] == 50360 && 
b[50361] == 50361 && 
b[50362] == 50362 && 
b[50363] == 50363 && 
b[50364] == 50364 && 
b[50365] == 50365 && 
b[50366] == 50366 && 
b[50367] == 50367 && 
b[50368] == 50368 && 
b[50369] == 50369 && 
b[50370] == 50370 && 
b[50371] == 50371 && 
b[50372] == 50372 && 
b[50373] == 50373 && 
b[50374] == 50374 && 
b[50375] == 50375 && 
b[50376] == 50376 && 
b[50377] == 50377 && 
b[50378] == 50378 && 
b[50379] == 50379 && 
b[50380] == 50380 && 
b[50381] == 50381 && 
b[50382] == 50382 && 
b[50383] == 50383 && 
b[50384] == 50384 && 
b[50385] == 50385 && 
b[50386] == 50386 && 
b[50387] == 50387 && 
b[50388] == 50388 && 
b[50389] == 50389 && 
b[50390] == 50390 && 
b[50391] == 50391 && 
b[50392] == 50392 && 
b[50393] == 50393 && 
b[50394] == 50394 && 
b[50395] == 50395 && 
b[50396] == 50396 && 
b[50397] == 50397 && 
b[50398] == 50398 && 
b[50399] == 50399 && 
b[50400] == 50400 && 
b[50401] == 50401 && 
b[50402] == 50402 && 
b[50403] == 50403 && 
b[50404] == 50404 && 
b[50405] == 50405 && 
b[50406] == 50406 && 
b[50407] == 50407 && 
b[50408] == 50408 && 
b[50409] == 50409 && 
b[50410] == 50410 && 
b[50411] == 50411 && 
b[50412] == 50412 && 
b[50413] == 50413 && 
b[50414] == 50414 && 
b[50415] == 50415 && 
b[50416] == 50416 && 
b[50417] == 50417 && 
b[50418] == 50418 && 
b[50419] == 50419 && 
b[50420] == 50420 && 
b[50421] == 50421 && 
b[50422] == 50422 && 
b[50423] == 50423 && 
b[50424] == 50424 && 
b[50425] == 50425 && 
b[50426] == 50426 && 
b[50427] == 50427 && 
b[50428] == 50428 && 
b[50429] == 50429 && 
b[50430] == 50430 && 
b[50431] == 50431 && 
b[50432] == 50432 && 
b[50433] == 50433 && 
b[50434] == 50434 && 
b[50435] == 50435 && 
b[50436] == 50436 && 
b[50437] == 50437 && 
b[50438] == 50438 && 
b[50439] == 50439 && 
b[50440] == 50440 && 
b[50441] == 50441 && 
b[50442] == 50442 && 
b[50443] == 50443 && 
b[50444] == 50444 && 
b[50445] == 50445 && 
b[50446] == 50446 && 
b[50447] == 50447 && 
b[50448] == 50448 && 
b[50449] == 50449 && 
b[50450] == 50450 && 
b[50451] == 50451 && 
b[50452] == 50452 && 
b[50453] == 50453 && 
b[50454] == 50454 && 
b[50455] == 50455 && 
b[50456] == 50456 && 
b[50457] == 50457 && 
b[50458] == 50458 && 
b[50459] == 50459 && 
b[50460] == 50460 && 
b[50461] == 50461 && 
b[50462] == 50462 && 
b[50463] == 50463 && 
b[50464] == 50464 && 
b[50465] == 50465 && 
b[50466] == 50466 && 
b[50467] == 50467 && 
b[50468] == 50468 && 
b[50469] == 50469 && 
b[50470] == 50470 && 
b[50471] == 50471 && 
b[50472] == 50472 && 
b[50473] == 50473 && 
b[50474] == 50474 && 
b[50475] == 50475 && 
b[50476] == 50476 && 
b[50477] == 50477 && 
b[50478] == 50478 && 
b[50479] == 50479 && 
b[50480] == 50480 && 
b[50481] == 50481 && 
b[50482] == 50482 && 
b[50483] == 50483 && 
b[50484] == 50484 && 
b[50485] == 50485 && 
b[50486] == 50486 && 
b[50487] == 50487 && 
b[50488] == 50488 && 
b[50489] == 50489 && 
b[50490] == 50490 && 
b[50491] == 50491 && 
b[50492] == 50492 && 
b[50493] == 50493 && 
b[50494] == 50494 && 
b[50495] == 50495 && 
b[50496] == 50496 && 
b[50497] == 50497 && 
b[50498] == 50498 && 
b[50499] == 50499 && 
b[50500] == 50500 && 
b[50501] == 50501 && 
b[50502] == 50502 && 
b[50503] == 50503 && 
b[50504] == 50504 && 
b[50505] == 50505 && 
b[50506] == 50506 && 
b[50507] == 50507 && 
b[50508] == 50508 && 
b[50509] == 50509 && 
b[50510] == 50510 && 
b[50511] == 50511 && 
b[50512] == 50512 && 
b[50513] == 50513 && 
b[50514] == 50514 && 
b[50515] == 50515 && 
b[50516] == 50516 && 
b[50517] == 50517 && 
b[50518] == 50518 && 
b[50519] == 50519 && 
b[50520] == 50520 && 
b[50521] == 50521 && 
b[50522] == 50522 && 
b[50523] == 50523 && 
b[50524] == 50524 && 
b[50525] == 50525 && 
b[50526] == 50526 && 
b[50527] == 50527 && 
b[50528] == 50528 && 
b[50529] == 50529 && 
b[50530] == 50530 && 
b[50531] == 50531 && 
b[50532] == 50532 && 
b[50533] == 50533 && 
b[50534] == 50534 && 
b[50535] == 50535 && 
b[50536] == 50536 && 
b[50537] == 50537 && 
b[50538] == 50538 && 
b[50539] == 50539 && 
b[50540] == 50540 && 
b[50541] == 50541 && 
b[50542] == 50542 && 
b[50543] == 50543 && 
b[50544] == 50544 && 
b[50545] == 50545 && 
b[50546] == 50546 && 
b[50547] == 50547 && 
b[50548] == 50548 && 
b[50549] == 50549 && 
b[50550] == 50550 && 
b[50551] == 50551 && 
b[50552] == 50552 && 
b[50553] == 50553 && 
b[50554] == 50554 && 
b[50555] == 50555 && 
b[50556] == 50556 && 
b[50557] == 50557 && 
b[50558] == 50558 && 
b[50559] == 50559 && 
b[50560] == 50560 && 
b[50561] == 50561 && 
b[50562] == 50562 && 
b[50563] == 50563 && 
b[50564] == 50564 && 
b[50565] == 50565 && 
b[50566] == 50566 && 
b[50567] == 50567 && 
b[50568] == 50568 && 
b[50569] == 50569 && 
b[50570] == 50570 && 
b[50571] == 50571 && 
b[50572] == 50572 && 
b[50573] == 50573 && 
b[50574] == 50574 && 
b[50575] == 50575 && 
b[50576] == 50576 && 
b[50577] == 50577 && 
b[50578] == 50578 && 
b[50579] == 50579 && 
b[50580] == 50580 && 
b[50581] == 50581 && 
b[50582] == 50582 && 
b[50583] == 50583 && 
b[50584] == 50584 && 
b[50585] == 50585 && 
b[50586] == 50586 && 
b[50587] == 50587 && 
b[50588] == 50588 && 
b[50589] == 50589 && 
b[50590] == 50590 && 
b[50591] == 50591 && 
b[50592] == 50592 && 
b[50593] == 50593 && 
b[50594] == 50594 && 
b[50595] == 50595 && 
b[50596] == 50596 && 
b[50597] == 50597 && 
b[50598] == 50598 && 
b[50599] == 50599 && 
b[50600] == 50600 && 
b[50601] == 50601 && 
b[50602] == 50602 && 
b[50603] == 50603 && 
b[50604] == 50604 && 
b[50605] == 50605 && 
b[50606] == 50606 && 
b[50607] == 50607 && 
b[50608] == 50608 && 
b[50609] == 50609 && 
b[50610] == 50610 && 
b[50611] == 50611 && 
b[50612] == 50612 && 
b[50613] == 50613 && 
b[50614] == 50614 && 
b[50615] == 50615 && 
b[50616] == 50616 && 
b[50617] == 50617 && 
b[50618] == 50618 && 
b[50619] == 50619 && 
b[50620] == 50620 && 
b[50621] == 50621 && 
b[50622] == 50622 && 
b[50623] == 50623 && 
b[50624] == 50624 && 
b[50625] == 50625 && 
b[50626] == 50626 && 
b[50627] == 50627 && 
b[50628] == 50628 && 
b[50629] == 50629 && 
b[50630] == 50630 && 
b[50631] == 50631 && 
b[50632] == 50632 && 
b[50633] == 50633 && 
b[50634] == 50634 && 
b[50635] == 50635 && 
b[50636] == 50636 && 
b[50637] == 50637 && 
b[50638] == 50638 && 
b[50639] == 50639 && 
b[50640] == 50640 && 
b[50641] == 50641 && 
b[50642] == 50642 && 
b[50643] == 50643 && 
b[50644] == 50644 && 
b[50645] == 50645 && 
b[50646] == 50646 && 
b[50647] == 50647 && 
b[50648] == 50648 && 
b[50649] == 50649 && 
b[50650] == 50650 && 
b[50651] == 50651 && 
b[50652] == 50652 && 
b[50653] == 50653 && 
b[50654] == 50654 && 
b[50655] == 50655 && 
b[50656] == 50656 && 
b[50657] == 50657 && 
b[50658] == 50658 && 
b[50659] == 50659 && 
b[50660] == 50660 && 
b[50661] == 50661 && 
b[50662] == 50662 && 
b[50663] == 50663 && 
b[50664] == 50664 && 
b[50665] == 50665 && 
b[50666] == 50666 && 
b[50667] == 50667 && 
b[50668] == 50668 && 
b[50669] == 50669 && 
b[50670] == 50670 && 
b[50671] == 50671 && 
b[50672] == 50672 && 
b[50673] == 50673 && 
b[50674] == 50674 && 
b[50675] == 50675 && 
b[50676] == 50676 && 
b[50677] == 50677 && 
b[50678] == 50678 && 
b[50679] == 50679 && 
b[50680] == 50680 && 
b[50681] == 50681 && 
b[50682] == 50682 && 
b[50683] == 50683 && 
b[50684] == 50684 && 
b[50685] == 50685 && 
b[50686] == 50686 && 
b[50687] == 50687 && 
b[50688] == 50688 && 
b[50689] == 50689 && 
b[50690] == 50690 && 
b[50691] == 50691 && 
b[50692] == 50692 && 
b[50693] == 50693 && 
b[50694] == 50694 && 
b[50695] == 50695 && 
b[50696] == 50696 && 
b[50697] == 50697 && 
b[50698] == 50698 && 
b[50699] == 50699 && 
b[50700] == 50700 && 
b[50701] == 50701 && 
b[50702] == 50702 && 
b[50703] == 50703 && 
b[50704] == 50704 && 
b[50705] == 50705 && 
b[50706] == 50706 && 
b[50707] == 50707 && 
b[50708] == 50708 && 
b[50709] == 50709 && 
b[50710] == 50710 && 
b[50711] == 50711 && 
b[50712] == 50712 && 
b[50713] == 50713 && 
b[50714] == 50714 && 
b[50715] == 50715 && 
b[50716] == 50716 && 
b[50717] == 50717 && 
b[50718] == 50718 && 
b[50719] == 50719 && 
b[50720] == 50720 && 
b[50721] == 50721 && 
b[50722] == 50722 && 
b[50723] == 50723 && 
b[50724] == 50724 && 
b[50725] == 50725 && 
b[50726] == 50726 && 
b[50727] == 50727 && 
b[50728] == 50728 && 
b[50729] == 50729 && 
b[50730] == 50730 && 
b[50731] == 50731 && 
b[50732] == 50732 && 
b[50733] == 50733 && 
b[50734] == 50734 && 
b[50735] == 50735 && 
b[50736] == 50736 && 
b[50737] == 50737 && 
b[50738] == 50738 && 
b[50739] == 50739 && 
b[50740] == 50740 && 
b[50741] == 50741 && 
b[50742] == 50742 && 
b[50743] == 50743 && 
b[50744] == 50744 && 
b[50745] == 50745 && 
b[50746] == 50746 && 
b[50747] == 50747 && 
b[50748] == 50748 && 
b[50749] == 50749 && 
b[50750] == 50750 && 
b[50751] == 50751 && 
b[50752] == 50752 && 
b[50753] == 50753 && 
b[50754] == 50754 && 
b[50755] == 50755 && 
b[50756] == 50756 && 
b[50757] == 50757 && 
b[50758] == 50758 && 
b[50759] == 50759 && 
b[50760] == 50760 && 
b[50761] == 50761 && 
b[50762] == 50762 && 
b[50763] == 50763 && 
b[50764] == 50764 && 
b[50765] == 50765 && 
b[50766] == 50766 && 
b[50767] == 50767 && 
b[50768] == 50768 && 
b[50769] == 50769 && 
b[50770] == 50770 && 
b[50771] == 50771 && 
b[50772] == 50772 && 
b[50773] == 50773 && 
b[50774] == 50774 && 
b[50775] == 50775 && 
b[50776] == 50776 && 
b[50777] == 50777 && 
b[50778] == 50778 && 
b[50779] == 50779 && 
b[50780] == 50780 && 
b[50781] == 50781 && 
b[50782] == 50782 && 
b[50783] == 50783 && 
b[50784] == 50784 && 
b[50785] == 50785 && 
b[50786] == 50786 && 
b[50787] == 50787 && 
b[50788] == 50788 && 
b[50789] == 50789 && 
b[50790] == 50790 && 
b[50791] == 50791 && 
b[50792] == 50792 && 
b[50793] == 50793 && 
b[50794] == 50794 && 
b[50795] == 50795 && 
b[50796] == 50796 && 
b[50797] == 50797 && 
b[50798] == 50798 && 
b[50799] == 50799 && 
b[50800] == 50800 && 
b[50801] == 50801 && 
b[50802] == 50802 && 
b[50803] == 50803 && 
b[50804] == 50804 && 
b[50805] == 50805 && 
b[50806] == 50806 && 
b[50807] == 50807 && 
b[50808] == 50808 && 
b[50809] == 50809 && 
b[50810] == 50810 && 
b[50811] == 50811 && 
b[50812] == 50812 && 
b[50813] == 50813 && 
b[50814] == 50814 && 
b[50815] == 50815 && 
b[50816] == 50816 && 
b[50817] == 50817 && 
b[50818] == 50818 && 
b[50819] == 50819 && 
b[50820] == 50820 && 
b[50821] == 50821 && 
b[50822] == 50822 && 
b[50823] == 50823 && 
b[50824] == 50824 && 
b[50825] == 50825 && 
b[50826] == 50826 && 
b[50827] == 50827 && 
b[50828] == 50828 && 
b[50829] == 50829 && 
b[50830] == 50830 && 
b[50831] == 50831 && 
b[50832] == 50832 && 
b[50833] == 50833 && 
b[50834] == 50834 && 
b[50835] == 50835 && 
b[50836] == 50836 && 
b[50837] == 50837 && 
b[50838] == 50838 && 
b[50839] == 50839 && 
b[50840] == 50840 && 
b[50841] == 50841 && 
b[50842] == 50842 && 
b[50843] == 50843 && 
b[50844] == 50844 && 
b[50845] == 50845 && 
b[50846] == 50846 && 
b[50847] == 50847 && 
b[50848] == 50848 && 
b[50849] == 50849 && 
b[50850] == 50850 && 
b[50851] == 50851 && 
b[50852] == 50852 && 
b[50853] == 50853 && 
b[50854] == 50854 && 
b[50855] == 50855 && 
b[50856] == 50856 && 
b[50857] == 50857 && 
b[50858] == 50858 && 
b[50859] == 50859 && 
b[50860] == 50860 && 
b[50861] == 50861 && 
b[50862] == 50862 && 
b[50863] == 50863 && 
b[50864] == 50864 && 
b[50865] == 50865 && 
b[50866] == 50866 && 
b[50867] == 50867 && 
b[50868] == 50868 && 
b[50869] == 50869 && 
b[50870] == 50870 && 
b[50871] == 50871 && 
b[50872] == 50872 && 
b[50873] == 50873 && 
b[50874] == 50874 && 
b[50875] == 50875 && 
b[50876] == 50876 && 
b[50877] == 50877 && 
b[50878] == 50878 && 
b[50879] == 50879 && 
b[50880] == 50880 && 
b[50881] == 50881 && 
b[50882] == 50882 && 
b[50883] == 50883 && 
b[50884] == 50884 && 
b[50885] == 50885 && 
b[50886] == 50886 && 
b[50887] == 50887 && 
b[50888] == 50888 && 
b[50889] == 50889 && 
b[50890] == 50890 && 
b[50891] == 50891 && 
b[50892] == 50892 && 
b[50893] == 50893 && 
b[50894] == 50894 && 
b[50895] == 50895 && 
b[50896] == 50896 && 
b[50897] == 50897 && 
b[50898] == 50898 && 
b[50899] == 50899 && 
b[50900] == 50900 && 
b[50901] == 50901 && 
b[50902] == 50902 && 
b[50903] == 50903 && 
b[50904] == 50904 && 
b[50905] == 50905 && 
b[50906] == 50906 && 
b[50907] == 50907 && 
b[50908] == 50908 && 
b[50909] == 50909 && 
b[50910] == 50910 && 
b[50911] == 50911 && 
b[50912] == 50912 && 
b[50913] == 50913 && 
b[50914] == 50914 && 
b[50915] == 50915 && 
b[50916] == 50916 && 
b[50917] == 50917 && 
b[50918] == 50918 && 
b[50919] == 50919 && 
b[50920] == 50920 && 
b[50921] == 50921 && 
b[50922] == 50922 && 
b[50923] == 50923 && 
b[50924] == 50924 && 
b[50925] == 50925 && 
b[50926] == 50926 && 
b[50927] == 50927 && 
b[50928] == 50928 && 
b[50929] == 50929 && 
b[50930] == 50930 && 
b[50931] == 50931 && 
b[50932] == 50932 && 
b[50933] == 50933 && 
b[50934] == 50934 && 
b[50935] == 50935 && 
b[50936] == 50936 && 
b[50937] == 50937 && 
b[50938] == 50938 && 
b[50939] == 50939 && 
b[50940] == 50940 && 
b[50941] == 50941 && 
b[50942] == 50942 && 
b[50943] == 50943 && 
b[50944] == 50944 && 
b[50945] == 50945 && 
b[50946] == 50946 && 
b[50947] == 50947 && 
b[50948] == 50948 && 
b[50949] == 50949 && 
b[50950] == 50950 && 
b[50951] == 50951 && 
b[50952] == 50952 && 
b[50953] == 50953 && 
b[50954] == 50954 && 
b[50955] == 50955 && 
b[50956] == 50956 && 
b[50957] == 50957 && 
b[50958] == 50958 && 
b[50959] == 50959 && 
b[50960] == 50960 && 
b[50961] == 50961 && 
b[50962] == 50962 && 
b[50963] == 50963 && 
b[50964] == 50964 && 
b[50965] == 50965 && 
b[50966] == 50966 && 
b[50967] == 50967 && 
b[50968] == 50968 && 
b[50969] == 50969 && 
b[50970] == 50970 && 
b[50971] == 50971 && 
b[50972] == 50972 && 
b[50973] == 50973 && 
b[50974] == 50974 && 
b[50975] == 50975 && 
b[50976] == 50976 && 
b[50977] == 50977 && 
b[50978] == 50978 && 
b[50979] == 50979 && 
b[50980] == 50980 && 
b[50981] == 50981 && 
b[50982] == 50982 && 
b[50983] == 50983 && 
b[50984] == 50984 && 
b[50985] == 50985 && 
b[50986] == 50986 && 
b[50987] == 50987 && 
b[50988] == 50988 && 
b[50989] == 50989 && 
b[50990] == 50990 && 
b[50991] == 50991 && 
b[50992] == 50992 && 
b[50993] == 50993 && 
b[50994] == 50994 && 
b[50995] == 50995 && 
b[50996] == 50996 && 
b[50997] == 50997 && 
b[50998] == 50998 && 
b[50999] == 50999 && 
b[51000] == 51000 && 
b[51001] == 51001 && 
b[51002] == 51002 && 
b[51003] == 51003 && 
b[51004] == 51004 && 
b[51005] == 51005 && 
b[51006] == 51006 && 
b[51007] == 51007 && 
b[51008] == 51008 && 
b[51009] == 51009 && 
b[51010] == 51010 && 
b[51011] == 51011 && 
b[51012] == 51012 && 
b[51013] == 51013 && 
b[51014] == 51014 && 
b[51015] == 51015 && 
b[51016] == 51016 && 
b[51017] == 51017 && 
b[51018] == 51018 && 
b[51019] == 51019 && 
b[51020] == 51020 && 
b[51021] == 51021 && 
b[51022] == 51022 && 
b[51023] == 51023 && 
b[51024] == 51024 && 
b[51025] == 51025 && 
b[51026] == 51026 && 
b[51027] == 51027 && 
b[51028] == 51028 && 
b[51029] == 51029 && 
b[51030] == 51030 && 
b[51031] == 51031 && 
b[51032] == 51032 && 
b[51033] == 51033 && 
b[51034] == 51034 && 
b[51035] == 51035 && 
b[51036] == 51036 && 
b[51037] == 51037 && 
b[51038] == 51038 && 
b[51039] == 51039 && 
b[51040] == 51040 && 
b[51041] == 51041 && 
b[51042] == 51042 && 
b[51043] == 51043 && 
b[51044] == 51044 && 
b[51045] == 51045 && 
b[51046] == 51046 && 
b[51047] == 51047 && 
b[51048] == 51048 && 
b[51049] == 51049 && 
b[51050] == 51050 && 
b[51051] == 51051 && 
b[51052] == 51052 && 
b[51053] == 51053 && 
b[51054] == 51054 && 
b[51055] == 51055 && 
b[51056] == 51056 && 
b[51057] == 51057 && 
b[51058] == 51058 && 
b[51059] == 51059 && 
b[51060] == 51060 && 
b[51061] == 51061 && 
b[51062] == 51062 && 
b[51063] == 51063 && 
b[51064] == 51064 && 
b[51065] == 51065 && 
b[51066] == 51066 && 
b[51067] == 51067 && 
b[51068] == 51068 && 
b[51069] == 51069 && 
b[51070] == 51070 && 
b[51071] == 51071 && 
b[51072] == 51072 && 
b[51073] == 51073 && 
b[51074] == 51074 && 
b[51075] == 51075 && 
b[51076] == 51076 && 
b[51077] == 51077 && 
b[51078] == 51078 && 
b[51079] == 51079 && 
b[51080] == 51080 && 
b[51081] == 51081 && 
b[51082] == 51082 && 
b[51083] == 51083 && 
b[51084] == 51084 && 
b[51085] == 51085 && 
b[51086] == 51086 && 
b[51087] == 51087 && 
b[51088] == 51088 && 
b[51089] == 51089 && 
b[51090] == 51090 && 
b[51091] == 51091 && 
b[51092] == 51092 && 
b[51093] == 51093 && 
b[51094] == 51094 && 
b[51095] == 51095 && 
b[51096] == 51096 && 
b[51097] == 51097 && 
b[51098] == 51098 && 
b[51099] == 51099 && 
b[51100] == 51100 && 
b[51101] == 51101 && 
b[51102] == 51102 && 
b[51103] == 51103 && 
b[51104] == 51104 && 
b[51105] == 51105 && 
b[51106] == 51106 && 
b[51107] == 51107 && 
b[51108] == 51108 && 
b[51109] == 51109 && 
b[51110] == 51110 && 
b[51111] == 51111 && 
b[51112] == 51112 && 
b[51113] == 51113 && 
b[51114] == 51114 && 
b[51115] == 51115 && 
b[51116] == 51116 && 
b[51117] == 51117 && 
b[51118] == 51118 && 
b[51119] == 51119 && 
b[51120] == 51120 && 
b[51121] == 51121 && 
b[51122] == 51122 && 
b[51123] == 51123 && 
b[51124] == 51124 && 
b[51125] == 51125 && 
b[51126] == 51126 && 
b[51127] == 51127 && 
b[51128] == 51128 && 
b[51129] == 51129 && 
b[51130] == 51130 && 
b[51131] == 51131 && 
b[51132] == 51132 && 
b[51133] == 51133 && 
b[51134] == 51134 && 
b[51135] == 51135 && 
b[51136] == 51136 && 
b[51137] == 51137 && 
b[51138] == 51138 && 
b[51139] == 51139 && 
b[51140] == 51140 && 
b[51141] == 51141 && 
b[51142] == 51142 && 
b[51143] == 51143 && 
b[51144] == 51144 && 
b[51145] == 51145 && 
b[51146] == 51146 && 
b[51147] == 51147 && 
b[51148] == 51148 && 
b[51149] == 51149 && 
b[51150] == 51150 && 
b[51151] == 51151 && 
b[51152] == 51152 && 
b[51153] == 51153 && 
b[51154] == 51154 && 
b[51155] == 51155 && 
b[51156] == 51156 && 
b[51157] == 51157 && 
b[51158] == 51158 && 
b[51159] == 51159 && 
b[51160] == 51160 && 
b[51161] == 51161 && 
b[51162] == 51162 && 
b[51163] == 51163 && 
b[51164] == 51164 && 
b[51165] == 51165 && 
b[51166] == 51166 && 
b[51167] == 51167 && 
b[51168] == 51168 && 
b[51169] == 51169 && 
b[51170] == 51170 && 
b[51171] == 51171 && 
b[51172] == 51172 && 
b[51173] == 51173 && 
b[51174] == 51174 && 
b[51175] == 51175 && 
b[51176] == 51176 && 
b[51177] == 51177 && 
b[51178] == 51178 && 
b[51179] == 51179 && 
b[51180] == 51180 && 
b[51181] == 51181 && 
b[51182] == 51182 && 
b[51183] == 51183 && 
b[51184] == 51184 && 
b[51185] == 51185 && 
b[51186] == 51186 && 
b[51187] == 51187 && 
b[51188] == 51188 && 
b[51189] == 51189 && 
b[51190] == 51190 && 
b[51191] == 51191 && 
b[51192] == 51192 && 
b[51193] == 51193 && 
b[51194] == 51194 && 
b[51195] == 51195 && 
b[51196] == 51196 && 
b[51197] == 51197 && 
b[51198] == 51198 && 
b[51199] == 51199 && 
b[51200] == 51200 && 
b[51201] == 51201 && 
b[51202] == 51202 && 
b[51203] == 51203 && 
b[51204] == 51204 && 
b[51205] == 51205 && 
b[51206] == 51206 && 
b[51207] == 51207 && 
b[51208] == 51208 && 
b[51209] == 51209 && 
b[51210] == 51210 && 
b[51211] == 51211 && 
b[51212] == 51212 && 
b[51213] == 51213 && 
b[51214] == 51214 && 
b[51215] == 51215 && 
b[51216] == 51216 && 
b[51217] == 51217 && 
b[51218] == 51218 && 
b[51219] == 51219 && 
b[51220] == 51220 && 
b[51221] == 51221 && 
b[51222] == 51222 && 
b[51223] == 51223 && 
b[51224] == 51224 && 
b[51225] == 51225 && 
b[51226] == 51226 && 
b[51227] == 51227 && 
b[51228] == 51228 && 
b[51229] == 51229 && 
b[51230] == 51230 && 
b[51231] == 51231 && 
b[51232] == 51232 && 
b[51233] == 51233 && 
b[51234] == 51234 && 
b[51235] == 51235 && 
b[51236] == 51236 && 
b[51237] == 51237 && 
b[51238] == 51238 && 
b[51239] == 51239 && 
b[51240] == 51240 && 
b[51241] == 51241 && 
b[51242] == 51242 && 
b[51243] == 51243 && 
b[51244] == 51244 && 
b[51245] == 51245 && 
b[51246] == 51246 && 
b[51247] == 51247 && 
b[51248] == 51248 && 
b[51249] == 51249 && 
b[51250] == 51250 && 
b[51251] == 51251 && 
b[51252] == 51252 && 
b[51253] == 51253 && 
b[51254] == 51254 && 
b[51255] == 51255 && 
b[51256] == 51256 && 
b[51257] == 51257 && 
b[51258] == 51258 && 
b[51259] == 51259 && 
b[51260] == 51260 && 
b[51261] == 51261 && 
b[51262] == 51262 && 
b[51263] == 51263 && 
b[51264] == 51264 && 
b[51265] == 51265 && 
b[51266] == 51266 && 
b[51267] == 51267 && 
b[51268] == 51268 && 
b[51269] == 51269 && 
b[51270] == 51270 && 
b[51271] == 51271 && 
b[51272] == 51272 && 
b[51273] == 51273 && 
b[51274] == 51274 && 
b[51275] == 51275 && 
b[51276] == 51276 && 
b[51277] == 51277 && 
b[51278] == 51278 && 
b[51279] == 51279 && 
b[51280] == 51280 && 
b[51281] == 51281 && 
b[51282] == 51282 && 
b[51283] == 51283 && 
b[51284] == 51284 && 
b[51285] == 51285 && 
b[51286] == 51286 && 
b[51287] == 51287 && 
b[51288] == 51288 && 
b[51289] == 51289 && 
b[51290] == 51290 && 
b[51291] == 51291 && 
b[51292] == 51292 && 
b[51293] == 51293 && 
b[51294] == 51294 && 
b[51295] == 51295 && 
b[51296] == 51296 && 
b[51297] == 51297 && 
b[51298] == 51298 && 
b[51299] == 51299 && 
b[51300] == 51300 && 
b[51301] == 51301 && 
b[51302] == 51302 && 
b[51303] == 51303 && 
b[51304] == 51304 && 
b[51305] == 51305 && 
b[51306] == 51306 && 
b[51307] == 51307 && 
b[51308] == 51308 && 
b[51309] == 51309 && 
b[51310] == 51310 && 
b[51311] == 51311 && 
b[51312] == 51312 && 
b[51313] == 51313 && 
b[51314] == 51314 && 
b[51315] == 51315 && 
b[51316] == 51316 && 
b[51317] == 51317 && 
b[51318] == 51318 && 
b[51319] == 51319 && 
b[51320] == 51320 && 
b[51321] == 51321 && 
b[51322] == 51322 && 
b[51323] == 51323 && 
b[51324] == 51324 && 
b[51325] == 51325 && 
b[51326] == 51326 && 
b[51327] == 51327 && 
b[51328] == 51328 && 
b[51329] == 51329 && 
b[51330] == 51330 && 
b[51331] == 51331 && 
b[51332] == 51332 && 
b[51333] == 51333 && 
b[51334] == 51334 && 
b[51335] == 51335 && 
b[51336] == 51336 && 
b[51337] == 51337 && 
b[51338] == 51338 && 
b[51339] == 51339 && 
b[51340] == 51340 && 
b[51341] == 51341 && 
b[51342] == 51342 && 
b[51343] == 51343 && 
b[51344] == 51344 && 
b[51345] == 51345 && 
b[51346] == 51346 && 
b[51347] == 51347 && 
b[51348] == 51348 && 
b[51349] == 51349 && 
b[51350] == 51350 && 
b[51351] == 51351 && 
b[51352] == 51352 && 
b[51353] == 51353 && 
b[51354] == 51354 && 
b[51355] == 51355 && 
b[51356] == 51356 && 
b[51357] == 51357 && 
b[51358] == 51358 && 
b[51359] == 51359 && 
b[51360] == 51360 && 
b[51361] == 51361 && 
b[51362] == 51362 && 
b[51363] == 51363 && 
b[51364] == 51364 && 
b[51365] == 51365 && 
b[51366] == 51366 && 
b[51367] == 51367 && 
b[51368] == 51368 && 
b[51369] == 51369 && 
b[51370] == 51370 && 
b[51371] == 51371 && 
b[51372] == 51372 && 
b[51373] == 51373 && 
b[51374] == 51374 && 
b[51375] == 51375 && 
b[51376] == 51376 && 
b[51377] == 51377 && 
b[51378] == 51378 && 
b[51379] == 51379 && 
b[51380] == 51380 && 
b[51381] == 51381 && 
b[51382] == 51382 && 
b[51383] == 51383 && 
b[51384] == 51384 && 
b[51385] == 51385 && 
b[51386] == 51386 && 
b[51387] == 51387 && 
b[51388] == 51388 && 
b[51389] == 51389 && 
b[51390] == 51390 && 
b[51391] == 51391 && 
b[51392] == 51392 && 
b[51393] == 51393 && 
b[51394] == 51394 && 
b[51395] == 51395 && 
b[51396] == 51396 && 
b[51397] == 51397 && 
b[51398] == 51398 && 
b[51399] == 51399 && 
b[51400] == 51400 && 
b[51401] == 51401 && 
b[51402] == 51402 && 
b[51403] == 51403 && 
b[51404] == 51404 && 
b[51405] == 51405 && 
b[51406] == 51406 && 
b[51407] == 51407 && 
b[51408] == 51408 && 
b[51409] == 51409 && 
b[51410] == 51410 && 
b[51411] == 51411 && 
b[51412] == 51412 && 
b[51413] == 51413 && 
b[51414] == 51414 && 
b[51415] == 51415 && 
b[51416] == 51416 && 
b[51417] == 51417 && 
b[51418] == 51418 && 
b[51419] == 51419 && 
b[51420] == 51420 && 
b[51421] == 51421 && 
b[51422] == 51422 && 
b[51423] == 51423 && 
b[51424] == 51424 && 
b[51425] == 51425 && 
b[51426] == 51426 && 
b[51427] == 51427 && 
b[51428] == 51428 && 
b[51429] == 51429 && 
b[51430] == 51430 && 
b[51431] == 51431 && 
b[51432] == 51432 && 
b[51433] == 51433 && 
b[51434] == 51434 && 
b[51435] == 51435 && 
b[51436] == 51436 && 
b[51437] == 51437 && 
b[51438] == 51438 && 
b[51439] == 51439 && 
b[51440] == 51440 && 
b[51441] == 51441 && 
b[51442] == 51442 && 
b[51443] == 51443 && 
b[51444] == 51444 && 
b[51445] == 51445 && 
b[51446] == 51446 && 
b[51447] == 51447 && 
b[51448] == 51448 && 
b[51449] == 51449 && 
b[51450] == 51450 && 
b[51451] == 51451 && 
b[51452] == 51452 && 
b[51453] == 51453 && 
b[51454] == 51454 && 
b[51455] == 51455 && 
b[51456] == 51456 && 
b[51457] == 51457 && 
b[51458] == 51458 && 
b[51459] == 51459 && 
b[51460] == 51460 && 
b[51461] == 51461 && 
b[51462] == 51462 && 
b[51463] == 51463 && 
b[51464] == 51464 && 
b[51465] == 51465 && 
b[51466] == 51466 && 
b[51467] == 51467 && 
b[51468] == 51468 && 
b[51469] == 51469 && 
b[51470] == 51470 && 
b[51471] == 51471 && 
b[51472] == 51472 && 
b[51473] == 51473 && 
b[51474] == 51474 && 
b[51475] == 51475 && 
b[51476] == 51476 && 
b[51477] == 51477 && 
b[51478] == 51478 && 
b[51479] == 51479 && 
b[51480] == 51480 && 
b[51481] == 51481 && 
b[51482] == 51482 && 
b[51483] == 51483 && 
b[51484] == 51484 && 
b[51485] == 51485 && 
b[51486] == 51486 && 
b[51487] == 51487 && 
b[51488] == 51488 && 
b[51489] == 51489 && 
b[51490] == 51490 && 
b[51491] == 51491 && 
b[51492] == 51492 && 
b[51493] == 51493 && 
b[51494] == 51494 && 
b[51495] == 51495 && 
b[51496] == 51496 && 
b[51497] == 51497 && 
b[51498] == 51498 && 
b[51499] == 51499 && 
b[51500] == 51500 && 
b[51501] == 51501 && 
b[51502] == 51502 && 
b[51503] == 51503 && 
b[51504] == 51504 && 
b[51505] == 51505 && 
b[51506] == 51506 && 
b[51507] == 51507 && 
b[51508] == 51508 && 
b[51509] == 51509 && 
b[51510] == 51510 && 
b[51511] == 51511 && 
b[51512] == 51512 && 
b[51513] == 51513 && 
b[51514] == 51514 && 
b[51515] == 51515 && 
b[51516] == 51516 && 
b[51517] == 51517 && 
b[51518] == 51518 && 
b[51519] == 51519 && 
b[51520] == 51520 && 
b[51521] == 51521 && 
b[51522] == 51522 && 
b[51523] == 51523 && 
b[51524] == 51524 && 
b[51525] == 51525 && 
b[51526] == 51526 && 
b[51527] == 51527 && 
b[51528] == 51528 && 
b[51529] == 51529 && 
b[51530] == 51530 && 
b[51531] == 51531 && 
b[51532] == 51532 && 
b[51533] == 51533 && 
b[51534] == 51534 && 
b[51535] == 51535 && 
b[51536] == 51536 && 
b[51537] == 51537 && 
b[51538] == 51538 && 
b[51539] == 51539 && 
b[51540] == 51540 && 
b[51541] == 51541 && 
b[51542] == 51542 && 
b[51543] == 51543 && 
b[51544] == 51544 && 
b[51545] == 51545 && 
b[51546] == 51546 && 
b[51547] == 51547 && 
b[51548] == 51548 && 
b[51549] == 51549 && 
b[51550] == 51550 && 
b[51551] == 51551 && 
b[51552] == 51552 && 
b[51553] == 51553 && 
b[51554] == 51554 && 
b[51555] == 51555 && 
b[51556] == 51556 && 
b[51557] == 51557 && 
b[51558] == 51558 && 
b[51559] == 51559 && 
b[51560] == 51560 && 
b[51561] == 51561 && 
b[51562] == 51562 && 
b[51563] == 51563 && 
b[51564] == 51564 && 
b[51565] == 51565 && 
b[51566] == 51566 && 
b[51567] == 51567 && 
b[51568] == 51568 && 
b[51569] == 51569 && 
b[51570] == 51570 && 
b[51571] == 51571 && 
b[51572] == 51572 && 
b[51573] == 51573 && 
b[51574] == 51574 && 
b[51575] == 51575 && 
b[51576] == 51576 && 
b[51577] == 51577 && 
b[51578] == 51578 && 
b[51579] == 51579 && 
b[51580] == 51580 && 
b[51581] == 51581 && 
b[51582] == 51582 && 
b[51583] == 51583 && 
b[51584] == 51584 && 
b[51585] == 51585 && 
b[51586] == 51586 && 
b[51587] == 51587 && 
b[51588] == 51588 && 
b[51589] == 51589 && 
b[51590] == 51590 && 
b[51591] == 51591 && 
b[51592] == 51592 && 
b[51593] == 51593 && 
b[51594] == 51594 && 
b[51595] == 51595 && 
b[51596] == 51596 && 
b[51597] == 51597 && 
b[51598] == 51598 && 
b[51599] == 51599 && 
b[51600] == 51600 && 
b[51601] == 51601 && 
b[51602] == 51602 && 
b[51603] == 51603 && 
b[51604] == 51604 && 
b[51605] == 51605 && 
b[51606] == 51606 && 
b[51607] == 51607 && 
b[51608] == 51608 && 
b[51609] == 51609 && 
b[51610] == 51610 && 
b[51611] == 51611 && 
b[51612] == 51612 && 
b[51613] == 51613 && 
b[51614] == 51614 && 
b[51615] == 51615 && 
b[51616] == 51616 && 
b[51617] == 51617 && 
b[51618] == 51618 && 
b[51619] == 51619 && 
b[51620] == 51620 && 
b[51621] == 51621 && 
b[51622] == 51622 && 
b[51623] == 51623 && 
b[51624] == 51624 && 
b[51625] == 51625 && 
b[51626] == 51626 && 
b[51627] == 51627 && 
b[51628] == 51628 && 
b[51629] == 51629 && 
b[51630] == 51630 && 
b[51631] == 51631 && 
b[51632] == 51632 && 
b[51633] == 51633 && 
b[51634] == 51634 && 
b[51635] == 51635 && 
b[51636] == 51636 && 
b[51637] == 51637 && 
b[51638] == 51638 && 
b[51639] == 51639 && 
b[51640] == 51640 && 
b[51641] == 51641 && 
b[51642] == 51642 && 
b[51643] == 51643 && 
b[51644] == 51644 && 
b[51645] == 51645 && 
b[51646] == 51646 && 
b[51647] == 51647 && 
b[51648] == 51648 && 
b[51649] == 51649 && 
b[51650] == 51650 && 
b[51651] == 51651 && 
b[51652] == 51652 && 
b[51653] == 51653 && 
b[51654] == 51654 && 
b[51655] == 51655 && 
b[51656] == 51656 && 
b[51657] == 51657 && 
b[51658] == 51658 && 
b[51659] == 51659 && 
b[51660] == 51660 && 
b[51661] == 51661 && 
b[51662] == 51662 && 
b[51663] == 51663 && 
b[51664] == 51664 && 
b[51665] == 51665 && 
b[51666] == 51666 && 
b[51667] == 51667 && 
b[51668] == 51668 && 
b[51669] == 51669 && 
b[51670] == 51670 && 
b[51671] == 51671 && 
b[51672] == 51672 && 
b[51673] == 51673 && 
b[51674] == 51674 && 
b[51675] == 51675 && 
b[51676] == 51676 && 
b[51677] == 51677 && 
b[51678] == 51678 && 
b[51679] == 51679 && 
b[51680] == 51680 && 
b[51681] == 51681 && 
b[51682] == 51682 && 
b[51683] == 51683 && 
b[51684] == 51684 && 
b[51685] == 51685 && 
b[51686] == 51686 && 
b[51687] == 51687 && 
b[51688] == 51688 && 
b[51689] == 51689 && 
b[51690] == 51690 && 
b[51691] == 51691 && 
b[51692] == 51692 && 
b[51693] == 51693 && 
b[51694] == 51694 && 
b[51695] == 51695 && 
b[51696] == 51696 && 
b[51697] == 51697 && 
b[51698] == 51698 && 
b[51699] == 51699 && 
b[51700] == 51700 && 
b[51701] == 51701 && 
b[51702] == 51702 && 
b[51703] == 51703 && 
b[51704] == 51704 && 
b[51705] == 51705 && 
b[51706] == 51706 && 
b[51707] == 51707 && 
b[51708] == 51708 && 
b[51709] == 51709 && 
b[51710] == 51710 && 
b[51711] == 51711 && 
b[51712] == 51712 && 
b[51713] == 51713 && 
b[51714] == 51714 && 
b[51715] == 51715 && 
b[51716] == 51716 && 
b[51717] == 51717 && 
b[51718] == 51718 && 
b[51719] == 51719 && 
b[51720] == 51720 && 
b[51721] == 51721 && 
b[51722] == 51722 && 
b[51723] == 51723 && 
b[51724] == 51724 && 
b[51725] == 51725 && 
b[51726] == 51726 && 
b[51727] == 51727 && 
b[51728] == 51728 && 
b[51729] == 51729 && 
b[51730] == 51730 && 
b[51731] == 51731 && 
b[51732] == 51732 && 
b[51733] == 51733 && 
b[51734] == 51734 && 
b[51735] == 51735 && 
b[51736] == 51736 && 
b[51737] == 51737 && 
b[51738] == 51738 && 
b[51739] == 51739 && 
b[51740] == 51740 && 
b[51741] == 51741 && 
b[51742] == 51742 && 
b[51743] == 51743 && 
b[51744] == 51744 && 
b[51745] == 51745 && 
b[51746] == 51746 && 
b[51747] == 51747 && 
b[51748] == 51748 && 
b[51749] == 51749 && 
b[51750] == 51750 && 
b[51751] == 51751 && 
b[51752] == 51752 && 
b[51753] == 51753 && 
b[51754] == 51754 && 
b[51755] == 51755 && 
b[51756] == 51756 && 
b[51757] == 51757 && 
b[51758] == 51758 && 
b[51759] == 51759 && 
b[51760] == 51760 && 
b[51761] == 51761 && 
b[51762] == 51762 && 
b[51763] == 51763 && 
b[51764] == 51764 && 
b[51765] == 51765 && 
b[51766] == 51766 && 
b[51767] == 51767 && 
b[51768] == 51768 && 
b[51769] == 51769 && 
b[51770] == 51770 && 
b[51771] == 51771 && 
b[51772] == 51772 && 
b[51773] == 51773 && 
b[51774] == 51774 && 
b[51775] == 51775 && 
b[51776] == 51776 && 
b[51777] == 51777 && 
b[51778] == 51778 && 
b[51779] == 51779 && 
b[51780] == 51780 && 
b[51781] == 51781 && 
b[51782] == 51782 && 
b[51783] == 51783 && 
b[51784] == 51784 && 
b[51785] == 51785 && 
b[51786] == 51786 && 
b[51787] == 51787 && 
b[51788] == 51788 && 
b[51789] == 51789 && 
b[51790] == 51790 && 
b[51791] == 51791 && 
b[51792] == 51792 && 
b[51793] == 51793 && 
b[51794] == 51794 && 
b[51795] == 51795 && 
b[51796] == 51796 && 
b[51797] == 51797 && 
b[51798] == 51798 && 
b[51799] == 51799 && 
b[51800] == 51800 && 
b[51801] == 51801 && 
b[51802] == 51802 && 
b[51803] == 51803 && 
b[51804] == 51804 && 
b[51805] == 51805 && 
b[51806] == 51806 && 
b[51807] == 51807 && 
b[51808] == 51808 && 
b[51809] == 51809 && 
b[51810] == 51810 && 
b[51811] == 51811 && 
b[51812] == 51812 && 
b[51813] == 51813 && 
b[51814] == 51814 && 
b[51815] == 51815 && 
b[51816] == 51816 && 
b[51817] == 51817 && 
b[51818] == 51818 && 
b[51819] == 51819 && 
b[51820] == 51820 && 
b[51821] == 51821 && 
b[51822] == 51822 && 
b[51823] == 51823 && 
b[51824] == 51824 && 
b[51825] == 51825 && 
b[51826] == 51826 && 
b[51827] == 51827 && 
b[51828] == 51828 && 
b[51829] == 51829 && 
b[51830] == 51830 && 
b[51831] == 51831 && 
b[51832] == 51832 && 
b[51833] == 51833 && 
b[51834] == 51834 && 
b[51835] == 51835 && 
b[51836] == 51836 && 
b[51837] == 51837 && 
b[51838] == 51838 && 
b[51839] == 51839 && 
b[51840] == 51840 && 
b[51841] == 51841 && 
b[51842] == 51842 && 
b[51843] == 51843 && 
b[51844] == 51844 && 
b[51845] == 51845 && 
b[51846] == 51846 && 
b[51847] == 51847 && 
b[51848] == 51848 && 
b[51849] == 51849 && 
b[51850] == 51850 && 
b[51851] == 51851 && 
b[51852] == 51852 && 
b[51853] == 51853 && 
b[51854] == 51854 && 
b[51855] == 51855 && 
b[51856] == 51856 && 
b[51857] == 51857 && 
b[51858] == 51858 && 
b[51859] == 51859 && 
b[51860] == 51860 && 
b[51861] == 51861 && 
b[51862] == 51862 && 
b[51863] == 51863 && 
b[51864] == 51864 && 
b[51865] == 51865 && 
b[51866] == 51866 && 
b[51867] == 51867 && 
b[51868] == 51868 && 
b[51869] == 51869 && 
b[51870] == 51870 && 
b[51871] == 51871 && 
b[51872] == 51872 && 
b[51873] == 51873 && 
b[51874] == 51874 && 
b[51875] == 51875 && 
b[51876] == 51876 && 
b[51877] == 51877 && 
b[51878] == 51878 && 
b[51879] == 51879 && 
b[51880] == 51880 && 
b[51881] == 51881 && 
b[51882] == 51882 && 
b[51883] == 51883 && 
b[51884] == 51884 && 
b[51885] == 51885 && 
b[51886] == 51886 && 
b[51887] == 51887 && 
b[51888] == 51888 && 
b[51889] == 51889 && 
b[51890] == 51890 && 
b[51891] == 51891 && 
b[51892] == 51892 && 
b[51893] == 51893 && 
b[51894] == 51894 && 
b[51895] == 51895 && 
b[51896] == 51896 && 
b[51897] == 51897 && 
b[51898] == 51898 && 
b[51899] == 51899 && 
b[51900] == 51900 && 
b[51901] == 51901 && 
b[51902] == 51902 && 
b[51903] == 51903 && 
b[51904] == 51904 && 
b[51905] == 51905 && 
b[51906] == 51906 && 
b[51907] == 51907 && 
b[51908] == 51908 && 
b[51909] == 51909 && 
b[51910] == 51910 && 
b[51911] == 51911 && 
b[51912] == 51912 && 
b[51913] == 51913 && 
b[51914] == 51914 && 
b[51915] == 51915 && 
b[51916] == 51916 && 
b[51917] == 51917 && 
b[51918] == 51918 && 
b[51919] == 51919 && 
b[51920] == 51920 && 
b[51921] == 51921 && 
b[51922] == 51922 && 
b[51923] == 51923 && 
b[51924] == 51924 && 
b[51925] == 51925 && 
b[51926] == 51926 && 
b[51927] == 51927 && 
b[51928] == 51928 && 
b[51929] == 51929 && 
b[51930] == 51930 && 
b[51931] == 51931 && 
b[51932] == 51932 && 
b[51933] == 51933 && 
b[51934] == 51934 && 
b[51935] == 51935 && 
b[51936] == 51936 && 
b[51937] == 51937 && 
b[51938] == 51938 && 
b[51939] == 51939 && 
b[51940] == 51940 && 
b[51941] == 51941 && 
b[51942] == 51942 && 
b[51943] == 51943 && 
b[51944] == 51944 && 
b[51945] == 51945 && 
b[51946] == 51946 && 
b[51947] == 51947 && 
b[51948] == 51948 && 
b[51949] == 51949 && 
b[51950] == 51950 && 
b[51951] == 51951 && 
b[51952] == 51952 && 
b[51953] == 51953 && 
b[51954] == 51954 && 
b[51955] == 51955 && 
b[51956] == 51956 && 
b[51957] == 51957 && 
b[51958] == 51958 && 
b[51959] == 51959 && 
b[51960] == 51960 && 
b[51961] == 51961 && 
b[51962] == 51962 && 
b[51963] == 51963 && 
b[51964] == 51964 && 
b[51965] == 51965 && 
b[51966] == 51966 && 
b[51967] == 51967 && 
b[51968] == 51968 && 
b[51969] == 51969 && 
b[51970] == 51970 && 
b[51971] == 51971 && 
b[51972] == 51972 && 
b[51973] == 51973 && 
b[51974] == 51974 && 
b[51975] == 51975 && 
b[51976] == 51976 && 
b[51977] == 51977 && 
b[51978] == 51978 && 
b[51979] == 51979 && 
b[51980] == 51980 && 
b[51981] == 51981 && 
b[51982] == 51982 && 
b[51983] == 51983 && 
b[51984] == 51984 && 
b[51985] == 51985 && 
b[51986] == 51986 && 
b[51987] == 51987 && 
b[51988] == 51988 && 
b[51989] == 51989 && 
b[51990] == 51990 && 
b[51991] == 51991 && 
b[51992] == 51992 && 
b[51993] == 51993 && 
b[51994] == 51994 && 
b[51995] == 51995 && 
b[51996] == 51996 && 
b[51997] == 51997 && 
b[51998] == 51998 && 
b[51999] == 51999 && 
b[52000] == 52000 && 
b[52001] == 52001 && 
b[52002] == 52002 && 
b[52003] == 52003 && 
b[52004] == 52004 && 
b[52005] == 52005 && 
b[52006] == 52006 && 
b[52007] == 52007 && 
b[52008] == 52008 && 
b[52009] == 52009 && 
b[52010] == 52010 && 
b[52011] == 52011 && 
b[52012] == 52012 && 
b[52013] == 52013 && 
b[52014] == 52014 && 
b[52015] == 52015 && 
b[52016] == 52016 && 
b[52017] == 52017 && 
b[52018] == 52018 && 
b[52019] == 52019 && 
b[52020] == 52020 && 
b[52021] == 52021 && 
b[52022] == 52022 && 
b[52023] == 52023 && 
b[52024] == 52024 && 
b[52025] == 52025 && 
b[52026] == 52026 && 
b[52027] == 52027 && 
b[52028] == 52028 && 
b[52029] == 52029 && 
b[52030] == 52030 && 
b[52031] == 52031 && 
b[52032] == 52032 && 
b[52033] == 52033 && 
b[52034] == 52034 && 
b[52035] == 52035 && 
b[52036] == 52036 && 
b[52037] == 52037 && 
b[52038] == 52038 && 
b[52039] == 52039 && 
b[52040] == 52040 && 
b[52041] == 52041 && 
b[52042] == 52042 && 
b[52043] == 52043 && 
b[52044] == 52044 && 
b[52045] == 52045 && 
b[52046] == 52046 && 
b[52047] == 52047 && 
b[52048] == 52048 && 
b[52049] == 52049 && 
b[52050] == 52050 && 
b[52051] == 52051 && 
b[52052] == 52052 && 
b[52053] == 52053 && 
b[52054] == 52054 && 
b[52055] == 52055 && 
b[52056] == 52056 && 
b[52057] == 52057 && 
b[52058] == 52058 && 
b[52059] == 52059 && 
b[52060] == 52060 && 
b[52061] == 52061 && 
b[52062] == 52062 && 
b[52063] == 52063 && 
b[52064] == 52064 && 
b[52065] == 52065 && 
b[52066] == 52066 && 
b[52067] == 52067 && 
b[52068] == 52068 && 
b[52069] == 52069 && 
b[52070] == 52070 && 
b[52071] == 52071 && 
b[52072] == 52072 && 
b[52073] == 52073 && 
b[52074] == 52074 && 
b[52075] == 52075 && 
b[52076] == 52076 && 
b[52077] == 52077 && 
b[52078] == 52078 && 
b[52079] == 52079 && 
b[52080] == 52080 && 
b[52081] == 52081 && 
b[52082] == 52082 && 
b[52083] == 52083 && 
b[52084] == 52084 && 
b[52085] == 52085 && 
b[52086] == 52086 && 
b[52087] == 52087 && 
b[52088] == 52088 && 
b[52089] == 52089 && 
b[52090] == 52090 && 
b[52091] == 52091 && 
b[52092] == 52092 && 
b[52093] == 52093 && 
b[52094] == 52094 && 
b[52095] == 52095 && 
b[52096] == 52096 && 
b[52097] == 52097 && 
b[52098] == 52098 && 
b[52099] == 52099 && 
b[52100] == 52100 && 
b[52101] == 52101 && 
b[52102] == 52102 && 
b[52103] == 52103 && 
b[52104] == 52104 && 
b[52105] == 52105 && 
b[52106] == 52106 && 
b[52107] == 52107 && 
b[52108] == 52108 && 
b[52109] == 52109 && 
b[52110] == 52110 && 
b[52111] == 52111 && 
b[52112] == 52112 && 
b[52113] == 52113 && 
b[52114] == 52114 && 
b[52115] == 52115 && 
b[52116] == 52116 && 
b[52117] == 52117 && 
b[52118] == 52118 && 
b[52119] == 52119 && 
b[52120] == 52120 && 
b[52121] == 52121 && 
b[52122] == 52122 && 
b[52123] == 52123 && 
b[52124] == 52124 && 
b[52125] == 52125 && 
b[52126] == 52126 && 
b[52127] == 52127 && 
b[52128] == 52128 && 
b[52129] == 52129 && 
b[52130] == 52130 && 
b[52131] == 52131 && 
b[52132] == 52132 && 
b[52133] == 52133 && 
b[52134] == 52134 && 
b[52135] == 52135 && 
b[52136] == 52136 && 
b[52137] == 52137 && 
b[52138] == 52138 && 
b[52139] == 52139 && 
b[52140] == 52140 && 
b[52141] == 52141 && 
b[52142] == 52142 && 
b[52143] == 52143 && 
b[52144] == 52144 && 
b[52145] == 52145 && 
b[52146] == 52146 && 
b[52147] == 52147 && 
b[52148] == 52148 && 
b[52149] == 52149 && 
b[52150] == 52150 && 
b[52151] == 52151 && 
b[52152] == 52152 && 
b[52153] == 52153 && 
b[52154] == 52154 && 
b[52155] == 52155 && 
b[52156] == 52156 && 
b[52157] == 52157 && 
b[52158] == 52158 && 
b[52159] == 52159 && 
b[52160] == 52160 && 
b[52161] == 52161 && 
b[52162] == 52162 && 
b[52163] == 52163 && 
b[52164] == 52164 && 
b[52165] == 52165 && 
b[52166] == 52166 && 
b[52167] == 52167 && 
b[52168] == 52168 && 
b[52169] == 52169 && 
b[52170] == 52170 && 
b[52171] == 52171 && 
b[52172] == 52172 && 
b[52173] == 52173 && 
b[52174] == 52174 && 
b[52175] == 52175 && 
b[52176] == 52176 && 
b[52177] == 52177 && 
b[52178] == 52178 && 
b[52179] == 52179 && 
b[52180] == 52180 && 
b[52181] == 52181 && 
b[52182] == 52182 && 
b[52183] == 52183 && 
b[52184] == 52184 && 
b[52185] == 52185 && 
b[52186] == 52186 && 
b[52187] == 52187 && 
b[52188] == 52188 && 
b[52189] == 52189 && 
b[52190] == 52190 && 
b[52191] == 52191 && 
b[52192] == 52192 && 
b[52193] == 52193 && 
b[52194] == 52194 && 
b[52195] == 52195 && 
b[52196] == 52196 && 
b[52197] == 52197 && 
b[52198] == 52198 && 
b[52199] == 52199 && 
b[52200] == 52200 && 
b[52201] == 52201 && 
b[52202] == 52202 && 
b[52203] == 52203 && 
b[52204] == 52204 && 
b[52205] == 52205 && 
b[52206] == 52206 && 
b[52207] == 52207 && 
b[52208] == 52208 && 
b[52209] == 52209 && 
b[52210] == 52210 && 
b[52211] == 52211 && 
b[52212] == 52212 && 
b[52213] == 52213 && 
b[52214] == 52214 && 
b[52215] == 52215 && 
b[52216] == 52216 && 
b[52217] == 52217 && 
b[52218] == 52218 && 
b[52219] == 52219 && 
b[52220] == 52220 && 
b[52221] == 52221 && 
b[52222] == 52222 && 
b[52223] == 52223 && 
b[52224] == 52224 && 
b[52225] == 52225 && 
b[52226] == 52226 && 
b[52227] == 52227 && 
b[52228] == 52228 && 
b[52229] == 52229 && 
b[52230] == 52230 && 
b[52231] == 52231 && 
b[52232] == 52232 && 
b[52233] == 52233 && 
b[52234] == 52234 && 
b[52235] == 52235 && 
b[52236] == 52236 && 
b[52237] == 52237 && 
b[52238] == 52238 && 
b[52239] == 52239 && 
b[52240] == 52240 && 
b[52241] == 52241 && 
b[52242] == 52242 && 
b[52243] == 52243 && 
b[52244] == 52244 && 
b[52245] == 52245 && 
b[52246] == 52246 && 
b[52247] == 52247 && 
b[52248] == 52248 && 
b[52249] == 52249 && 
b[52250] == 52250 && 
b[52251] == 52251 && 
b[52252] == 52252 && 
b[52253] == 52253 && 
b[52254] == 52254 && 
b[52255] == 52255 && 
b[52256] == 52256 && 
b[52257] == 52257 && 
b[52258] == 52258 && 
b[52259] == 52259 && 
b[52260] == 52260 && 
b[52261] == 52261 && 
b[52262] == 52262 && 
b[52263] == 52263 && 
b[52264] == 52264 && 
b[52265] == 52265 && 
b[52266] == 52266 && 
b[52267] == 52267 && 
b[52268] == 52268 && 
b[52269] == 52269 && 
b[52270] == 52270 && 
b[52271] == 52271 && 
b[52272] == 52272 && 
b[52273] == 52273 && 
b[52274] == 52274 && 
b[52275] == 52275 && 
b[52276] == 52276 && 
b[52277] == 52277 && 
b[52278] == 52278 && 
b[52279] == 52279 && 
b[52280] == 52280 && 
b[52281] == 52281 && 
b[52282] == 52282 && 
b[52283] == 52283 && 
b[52284] == 52284 && 
b[52285] == 52285 && 
b[52286] == 52286 && 
b[52287] == 52287 && 
b[52288] == 52288 && 
b[52289] == 52289 && 
b[52290] == 52290 && 
b[52291] == 52291 && 
b[52292] == 52292 && 
b[52293] == 52293 && 
b[52294] == 52294 && 
b[52295] == 52295 && 
b[52296] == 52296 && 
b[52297] == 52297 && 
b[52298] == 52298 && 
b[52299] == 52299 && 
b[52300] == 52300 && 
b[52301] == 52301 && 
b[52302] == 52302 && 
b[52303] == 52303 && 
b[52304] == 52304 && 
b[52305] == 52305 && 
b[52306] == 52306 && 
b[52307] == 52307 && 
b[52308] == 52308 && 
b[52309] == 52309 && 
b[52310] == 52310 && 
b[52311] == 52311 && 
b[52312] == 52312 && 
b[52313] == 52313 && 
b[52314] == 52314 && 
b[52315] == 52315 && 
b[52316] == 52316 && 
b[52317] == 52317 && 
b[52318] == 52318 && 
b[52319] == 52319 && 
b[52320] == 52320 && 
b[52321] == 52321 && 
b[52322] == 52322 && 
b[52323] == 52323 && 
b[52324] == 52324 && 
b[52325] == 52325 && 
b[52326] == 52326 && 
b[52327] == 52327 && 
b[52328] == 52328 && 
b[52329] == 52329 && 
b[52330] == 52330 && 
b[52331] == 52331 && 
b[52332] == 52332 && 
b[52333] == 52333 && 
b[52334] == 52334 && 
b[52335] == 52335 && 
b[52336] == 52336 && 
b[52337] == 52337 && 
b[52338] == 52338 && 
b[52339] == 52339 && 
b[52340] == 52340 && 
b[52341] == 52341 && 
b[52342] == 52342 && 
b[52343] == 52343 && 
b[52344] == 52344 && 
b[52345] == 52345 && 
b[52346] == 52346 && 
b[52347] == 52347 && 
b[52348] == 52348 && 
b[52349] == 52349 && 
b[52350] == 52350 && 
b[52351] == 52351 && 
b[52352] == 52352 && 
b[52353] == 52353 && 
b[52354] == 52354 && 
b[52355] == 52355 && 
b[52356] == 52356 && 
b[52357] == 52357 && 
b[52358] == 52358 && 
b[52359] == 52359 && 
b[52360] == 52360 && 
b[52361] == 52361 && 
b[52362] == 52362 && 
b[52363] == 52363 && 
b[52364] == 52364 && 
b[52365] == 52365 && 
b[52366] == 52366 && 
b[52367] == 52367 && 
b[52368] == 52368 && 
b[52369] == 52369 && 
b[52370] == 52370 && 
b[52371] == 52371 && 
b[52372] == 52372 && 
b[52373] == 52373 && 
b[52374] == 52374 && 
b[52375] == 52375 && 
b[52376] == 52376 && 
b[52377] == 52377 && 
b[52378] == 52378 && 
b[52379] == 52379 && 
b[52380] == 52380 && 
b[52381] == 52381 && 
b[52382] == 52382 && 
b[52383] == 52383 && 
b[52384] == 52384 && 
b[52385] == 52385 && 
b[52386] == 52386 && 
b[52387] == 52387 && 
b[52388] == 52388 && 
b[52389] == 52389 && 
b[52390] == 52390 && 
b[52391] == 52391 && 
b[52392] == 52392 && 
b[52393] == 52393 && 
b[52394] == 52394 && 
b[52395] == 52395 && 
b[52396] == 52396 && 
b[52397] == 52397 && 
b[52398] == 52398 && 
b[52399] == 52399 && 
b[52400] == 52400 && 
b[52401] == 52401 && 
b[52402] == 52402 && 
b[52403] == 52403 && 
b[52404] == 52404 && 
b[52405] == 52405 && 
b[52406] == 52406 && 
b[52407] == 52407 && 
b[52408] == 52408 && 
b[52409] == 52409 && 
b[52410] == 52410 && 
b[52411] == 52411 && 
b[52412] == 52412 && 
b[52413] == 52413 && 
b[52414] == 52414 && 
b[52415] == 52415 && 
b[52416] == 52416 && 
b[52417] == 52417 && 
b[52418] == 52418 && 
b[52419] == 52419 && 
b[52420] == 52420 && 
b[52421] == 52421 && 
b[52422] == 52422 && 
b[52423] == 52423 && 
b[52424] == 52424 && 
b[52425] == 52425 && 
b[52426] == 52426 && 
b[52427] == 52427 && 
b[52428] == 52428 && 
b[52429] == 52429 && 
b[52430] == 52430 && 
b[52431] == 52431 && 
b[52432] == 52432 && 
b[52433] == 52433 && 
b[52434] == 52434 && 
b[52435] == 52435 && 
b[52436] == 52436 && 
b[52437] == 52437 && 
b[52438] == 52438 && 
b[52439] == 52439 && 
b[52440] == 52440 && 
b[52441] == 52441 && 
b[52442] == 52442 && 
b[52443] == 52443 && 
b[52444] == 52444 && 
b[52445] == 52445 && 
b[52446] == 52446 && 
b[52447] == 52447 && 
b[52448] == 52448 && 
b[52449] == 52449 && 
b[52450] == 52450 && 
b[52451] == 52451 && 
b[52452] == 52452 && 
b[52453] == 52453 && 
b[52454] == 52454 && 
b[52455] == 52455 && 
b[52456] == 52456 && 
b[52457] == 52457 && 
b[52458] == 52458 && 
b[52459] == 52459 && 
b[52460] == 52460 && 
b[52461] == 52461 && 
b[52462] == 52462 && 
b[52463] == 52463 && 
b[52464] == 52464 && 
b[52465] == 52465 && 
b[52466] == 52466 && 
b[52467] == 52467 && 
b[52468] == 52468 && 
b[52469] == 52469 && 
b[52470] == 52470 && 
b[52471] == 52471 && 
b[52472] == 52472 && 
b[52473] == 52473 && 
b[52474] == 52474 && 
b[52475] == 52475 && 
b[52476] == 52476 && 
b[52477] == 52477 && 
b[52478] == 52478 && 
b[52479] == 52479 && 
b[52480] == 52480 && 
b[52481] == 52481 && 
b[52482] == 52482 && 
b[52483] == 52483 && 
b[52484] == 52484 && 
b[52485] == 52485 && 
b[52486] == 52486 && 
b[52487] == 52487 && 
b[52488] == 52488 && 
b[52489] == 52489 && 
b[52490] == 52490 && 
b[52491] == 52491 && 
b[52492] == 52492 && 
b[52493] == 52493 && 
b[52494] == 52494 && 
b[52495] == 52495 && 
b[52496] == 52496 && 
b[52497] == 52497 && 
b[52498] == 52498 && 
b[52499] == 52499 && 
b[52500] == 52500 && 
b[52501] == 52501 && 
b[52502] == 52502 && 
b[52503] == 52503 && 
b[52504] == 52504 && 
b[52505] == 52505 && 
b[52506] == 52506 && 
b[52507] == 52507 && 
b[52508] == 52508 && 
b[52509] == 52509 && 
b[52510] == 52510 && 
b[52511] == 52511 && 
b[52512] == 52512 && 
b[52513] == 52513 && 
b[52514] == 52514 && 
b[52515] == 52515 && 
b[52516] == 52516 && 
b[52517] == 52517 && 
b[52518] == 52518 && 
b[52519] == 52519 && 
b[52520] == 52520 && 
b[52521] == 52521 && 
b[52522] == 52522 && 
b[52523] == 52523 && 
b[52524] == 52524 && 
b[52525] == 52525 && 
b[52526] == 52526 && 
b[52527] == 52527 && 
b[52528] == 52528 && 
b[52529] == 52529 && 
b[52530] == 52530 && 
b[52531] == 52531 && 
b[52532] == 52532 && 
b[52533] == 52533 && 
b[52534] == 52534 && 
b[52535] == 52535 && 
b[52536] == 52536 && 
b[52537] == 52537 && 
b[52538] == 52538 && 
b[52539] == 52539 && 
b[52540] == 52540 && 
b[52541] == 52541 && 
b[52542] == 52542 && 
b[52543] == 52543 && 
b[52544] == 52544 && 
b[52545] == 52545 && 
b[52546] == 52546 && 
b[52547] == 52547 && 
b[52548] == 52548 && 
b[52549] == 52549 && 
b[52550] == 52550 && 
b[52551] == 52551 && 
b[52552] == 52552 && 
b[52553] == 52553 && 
b[52554] == 52554 && 
b[52555] == 52555 && 
b[52556] == 52556 && 
b[52557] == 52557 && 
b[52558] == 52558 && 
b[52559] == 52559 && 
b[52560] == 52560 && 
b[52561] == 52561 && 
b[52562] == 52562 && 
b[52563] == 52563 && 
b[52564] == 52564 && 
b[52565] == 52565 && 
b[52566] == 52566 && 
b[52567] == 52567 && 
b[52568] == 52568 && 
b[52569] == 52569 && 
b[52570] == 52570 && 
b[52571] == 52571 && 
b[52572] == 52572 && 
b[52573] == 52573 && 
b[52574] == 52574 && 
b[52575] == 52575 && 
b[52576] == 52576 && 
b[52577] == 52577 && 
b[52578] == 52578 && 
b[52579] == 52579 && 
b[52580] == 52580 && 
b[52581] == 52581 && 
b[52582] == 52582 && 
b[52583] == 52583 && 
b[52584] == 52584 && 
b[52585] == 52585 && 
b[52586] == 52586 && 
b[52587] == 52587 && 
b[52588] == 52588 && 
b[52589] == 52589 && 
b[52590] == 52590 && 
b[52591] == 52591 && 
b[52592] == 52592 && 
b[52593] == 52593 && 
b[52594] == 52594 && 
b[52595] == 52595 && 
b[52596] == 52596 && 
b[52597] == 52597 && 
b[52598] == 52598 && 
b[52599] == 52599 && 
b[52600] == 52600 && 
b[52601] == 52601 && 
b[52602] == 52602 && 
b[52603] == 52603 && 
b[52604] == 52604 && 
b[52605] == 52605 && 
b[52606] == 52606 && 
b[52607] == 52607 && 
b[52608] == 52608 && 
b[52609] == 52609 && 
b[52610] == 52610 && 
b[52611] == 52611 && 
b[52612] == 52612 && 
b[52613] == 52613 && 
b[52614] == 52614 && 
b[52615] == 52615 && 
b[52616] == 52616 && 
b[52617] == 52617 && 
b[52618] == 52618 && 
b[52619] == 52619 && 
b[52620] == 52620 && 
b[52621] == 52621 && 
b[52622] == 52622 && 
b[52623] == 52623 && 
b[52624] == 52624 && 
b[52625] == 52625 && 
b[52626] == 52626 && 
b[52627] == 52627 && 
b[52628] == 52628 && 
b[52629] == 52629 && 
b[52630] == 52630 && 
b[52631] == 52631 && 
b[52632] == 52632 && 
b[52633] == 52633 && 
b[52634] == 52634 && 
b[52635] == 52635 && 
b[52636] == 52636 && 
b[52637] == 52637 && 
b[52638] == 52638 && 
b[52639] == 52639 && 
b[52640] == 52640 && 
b[52641] == 52641 && 
b[52642] == 52642 && 
b[52643] == 52643 && 
b[52644] == 52644 && 
b[52645] == 52645 && 
b[52646] == 52646 && 
b[52647] == 52647 && 
b[52648] == 52648 && 
b[52649] == 52649 && 
b[52650] == 52650 && 
b[52651] == 52651 && 
b[52652] == 52652 && 
b[52653] == 52653 && 
b[52654] == 52654 && 
b[52655] == 52655 && 
b[52656] == 52656 && 
b[52657] == 52657 && 
b[52658] == 52658 && 
b[52659] == 52659 && 
b[52660] == 52660 && 
b[52661] == 52661 && 
b[52662] == 52662 && 
b[52663] == 52663 && 
b[52664] == 52664 && 
b[52665] == 52665 && 
b[52666] == 52666 && 
b[52667] == 52667 && 
b[52668] == 52668 && 
b[52669] == 52669 && 
b[52670] == 52670 && 
b[52671] == 52671 && 
b[52672] == 52672 && 
b[52673] == 52673 && 
b[52674] == 52674 && 
b[52675] == 52675 && 
b[52676] == 52676 && 
b[52677] == 52677 && 
b[52678] == 52678 && 
b[52679] == 52679 && 
b[52680] == 52680 && 
b[52681] == 52681 && 
b[52682] == 52682 && 
b[52683] == 52683 && 
b[52684] == 52684 && 
b[52685] == 52685 && 
b[52686] == 52686 && 
b[52687] == 52687 && 
b[52688] == 52688 && 
b[52689] == 52689 && 
b[52690] == 52690 && 
b[52691] == 52691 && 
b[52692] == 52692 && 
b[52693] == 52693 && 
b[52694] == 52694 && 
b[52695] == 52695 && 
b[52696] == 52696 && 
b[52697] == 52697 && 
b[52698] == 52698 && 
b[52699] == 52699 && 
b[52700] == 52700 && 
b[52701] == 52701 && 
b[52702] == 52702 && 
b[52703] == 52703 && 
b[52704] == 52704 && 
b[52705] == 52705 && 
b[52706] == 52706 && 
b[52707] == 52707 && 
b[52708] == 52708 && 
b[52709] == 52709 && 
b[52710] == 52710 && 
b[52711] == 52711 && 
b[52712] == 52712 && 
b[52713] == 52713 && 
b[52714] == 52714 && 
b[52715] == 52715 && 
b[52716] == 52716 && 
b[52717] == 52717 && 
b[52718] == 52718 && 
b[52719] == 52719 && 
b[52720] == 52720 && 
b[52721] == 52721 && 
b[52722] == 52722 && 
b[52723] == 52723 && 
b[52724] == 52724 && 
b[52725] == 52725 && 
b[52726] == 52726 && 
b[52727] == 52727 && 
b[52728] == 52728 && 
b[52729] == 52729 && 
b[52730] == 52730 && 
b[52731] == 52731 && 
b[52732] == 52732 && 
b[52733] == 52733 && 
b[52734] == 52734 && 
b[52735] == 52735 && 
b[52736] == 52736 && 
b[52737] == 52737 && 
b[52738] == 52738 && 
b[52739] == 52739 && 
b[52740] == 52740 && 
b[52741] == 52741 && 
b[52742] == 52742 && 
b[52743] == 52743 && 
b[52744] == 52744 && 
b[52745] == 52745 && 
b[52746] == 52746 && 
b[52747] == 52747 && 
b[52748] == 52748 && 
b[52749] == 52749 && 
b[52750] == 52750 && 
b[52751] == 52751 && 
b[52752] == 52752 && 
b[52753] == 52753 && 
b[52754] == 52754 && 
b[52755] == 52755 && 
b[52756] == 52756 && 
b[52757] == 52757 && 
b[52758] == 52758 && 
b[52759] == 52759 && 
b[52760] == 52760 && 
b[52761] == 52761 && 
b[52762] == 52762 && 
b[52763] == 52763 && 
b[52764] == 52764 && 
b[52765] == 52765 && 
b[52766] == 52766 && 
b[52767] == 52767 && 
b[52768] == 52768 && 
b[52769] == 52769 && 
b[52770] == 52770 && 
b[52771] == 52771 && 
b[52772] == 52772 && 
b[52773] == 52773 && 
b[52774] == 52774 && 
b[52775] == 52775 && 
b[52776] == 52776 && 
b[52777] == 52777 && 
b[52778] == 52778 && 
b[52779] == 52779 && 
b[52780] == 52780 && 
b[52781] == 52781 && 
b[52782] == 52782 && 
b[52783] == 52783 && 
b[52784] == 52784 && 
b[52785] == 52785 && 
b[52786] == 52786 && 
b[52787] == 52787 && 
b[52788] == 52788 && 
b[52789] == 52789 && 
b[52790] == 52790 && 
b[52791] == 52791 && 
b[52792] == 52792 && 
b[52793] == 52793 && 
b[52794] == 52794 && 
b[52795] == 52795 && 
b[52796] == 52796 && 
b[52797] == 52797 && 
b[52798] == 52798 && 
b[52799] == 52799 && 
b[52800] == 52800 && 
b[52801] == 52801 && 
b[52802] == 52802 && 
b[52803] == 52803 && 
b[52804] == 52804 && 
b[52805] == 52805 && 
b[52806] == 52806 && 
b[52807] == 52807 && 
b[52808] == 52808 && 
b[52809] == 52809 && 
b[52810] == 52810 && 
b[52811] == 52811 && 
b[52812] == 52812 && 
b[52813] == 52813 && 
b[52814] == 52814 && 
b[52815] == 52815 && 
b[52816] == 52816 && 
b[52817] == 52817 && 
b[52818] == 52818 && 
b[52819] == 52819 && 
b[52820] == 52820 && 
b[52821] == 52821 && 
b[52822] == 52822 && 
b[52823] == 52823 && 
b[52824] == 52824 && 
b[52825] == 52825 && 
b[52826] == 52826 && 
b[52827] == 52827 && 
b[52828] == 52828 && 
b[52829] == 52829 && 
b[52830] == 52830 && 
b[52831] == 52831 && 
b[52832] == 52832 && 
b[52833] == 52833 && 
b[52834] == 52834 && 
b[52835] == 52835 && 
b[52836] == 52836 && 
b[52837] == 52837 && 
b[52838] == 52838 && 
b[52839] == 52839 && 
b[52840] == 52840 && 
b[52841] == 52841 && 
b[52842] == 52842 && 
b[52843] == 52843 && 
b[52844] == 52844 && 
b[52845] == 52845 && 
b[52846] == 52846 && 
b[52847] == 52847 && 
b[52848] == 52848 && 
b[52849] == 52849 && 
b[52850] == 52850 && 
b[52851] == 52851 && 
b[52852] == 52852 && 
b[52853] == 52853 && 
b[52854] == 52854 && 
b[52855] == 52855 && 
b[52856] == 52856 && 
b[52857] == 52857 && 
b[52858] == 52858 && 
b[52859] == 52859 && 
b[52860] == 52860 && 
b[52861] == 52861 && 
b[52862] == 52862 && 
b[52863] == 52863 && 
b[52864] == 52864 && 
b[52865] == 52865 && 
b[52866] == 52866 && 
b[52867] == 52867 && 
b[52868] == 52868 && 
b[52869] == 52869 && 
b[52870] == 52870 && 
b[52871] == 52871 && 
b[52872] == 52872 && 
b[52873] == 52873 && 
b[52874] == 52874 && 
b[52875] == 52875 && 
b[52876] == 52876 && 
b[52877] == 52877 && 
b[52878] == 52878 && 
b[52879] == 52879 && 
b[52880] == 52880 && 
b[52881] == 52881 && 
b[52882] == 52882 && 
b[52883] == 52883 && 
b[52884] == 52884 && 
b[52885] == 52885 && 
b[52886] == 52886 && 
b[52887] == 52887 && 
b[52888] == 52888 && 
b[52889] == 52889 && 
b[52890] == 52890 && 
b[52891] == 52891 && 
b[52892] == 52892 && 
b[52893] == 52893 && 
b[52894] == 52894 && 
b[52895] == 52895 && 
b[52896] == 52896 && 
b[52897] == 52897 && 
b[52898] == 52898 && 
b[52899] == 52899 && 
b[52900] == 52900 && 
b[52901] == 52901 && 
b[52902] == 52902 && 
b[52903] == 52903 && 
b[52904] == 52904 && 
b[52905] == 52905 && 
b[52906] == 52906 && 
b[52907] == 52907 && 
b[52908] == 52908 && 
b[52909] == 52909 && 
b[52910] == 52910 && 
b[52911] == 52911 && 
b[52912] == 52912 && 
b[52913] == 52913 && 
b[52914] == 52914 && 
b[52915] == 52915 && 
b[52916] == 52916 && 
b[52917] == 52917 && 
b[52918] == 52918 && 
b[52919] == 52919 && 
b[52920] == 52920 && 
b[52921] == 52921 && 
b[52922] == 52922 && 
b[52923] == 52923 && 
b[52924] == 52924 && 
b[52925] == 52925 && 
b[52926] == 52926 && 
b[52927] == 52927 && 
b[52928] == 52928 && 
b[52929] == 52929 && 
b[52930] == 52930 && 
b[52931] == 52931 && 
b[52932] == 52932 && 
b[52933] == 52933 && 
b[52934] == 52934 && 
b[52935] == 52935 && 
b[52936] == 52936 && 
b[52937] == 52937 && 
b[52938] == 52938 && 
b[52939] == 52939 && 
b[52940] == 52940 && 
b[52941] == 52941 && 
b[52942] == 52942 && 
b[52943] == 52943 && 
b[52944] == 52944 && 
b[52945] == 52945 && 
b[52946] == 52946 && 
b[52947] == 52947 && 
b[52948] == 52948 && 
b[52949] == 52949 && 
b[52950] == 52950 && 
b[52951] == 52951 && 
b[52952] == 52952 && 
b[52953] == 52953 && 
b[52954] == 52954 && 
b[52955] == 52955 && 
b[52956] == 52956 && 
b[52957] == 52957 && 
b[52958] == 52958 && 
b[52959] == 52959 && 
b[52960] == 52960 && 
b[52961] == 52961 && 
b[52962] == 52962 && 
b[52963] == 52963 && 
b[52964] == 52964 && 
b[52965] == 52965 && 
b[52966] == 52966 && 
b[52967] == 52967 && 
b[52968] == 52968 && 
b[52969] == 52969 && 
b[52970] == 52970 && 
b[52971] == 52971 && 
b[52972] == 52972 && 
b[52973] == 52973 && 
b[52974] == 52974 && 
b[52975] == 52975 && 
b[52976] == 52976 && 
b[52977] == 52977 && 
b[52978] == 52978 && 
b[52979] == 52979 && 
b[52980] == 52980 && 
b[52981] == 52981 && 
b[52982] == 52982 && 
b[52983] == 52983 && 
b[52984] == 52984 && 
b[52985] == 52985 && 
b[52986] == 52986 && 
b[52987] == 52987 && 
b[52988] == 52988 && 
b[52989] == 52989 && 
b[52990] == 52990 && 
b[52991] == 52991 && 
b[52992] == 52992 && 
b[52993] == 52993 && 
b[52994] == 52994 && 
b[52995] == 52995 && 
b[52996] == 52996 && 
b[52997] == 52997 && 
b[52998] == 52998 && 
b[52999] == 52999 && 
b[53000] == 53000 && 
b[53001] == 53001 && 
b[53002] == 53002 && 
b[53003] == 53003 && 
b[53004] == 53004 && 
b[53005] == 53005 && 
b[53006] == 53006 && 
b[53007] == 53007 && 
b[53008] == 53008 && 
b[53009] == 53009 && 
b[53010] == 53010 && 
b[53011] == 53011 && 
b[53012] == 53012 && 
b[53013] == 53013 && 
b[53014] == 53014 && 
b[53015] == 53015 && 
b[53016] == 53016 && 
b[53017] == 53017 && 
b[53018] == 53018 && 
b[53019] == 53019 && 
b[53020] == 53020 && 
b[53021] == 53021 && 
b[53022] == 53022 && 
b[53023] == 53023 && 
b[53024] == 53024 && 
b[53025] == 53025 && 
b[53026] == 53026 && 
b[53027] == 53027 && 
b[53028] == 53028 && 
b[53029] == 53029 && 
b[53030] == 53030 && 
b[53031] == 53031 && 
b[53032] == 53032 && 
b[53033] == 53033 && 
b[53034] == 53034 && 
b[53035] == 53035 && 
b[53036] == 53036 && 
b[53037] == 53037 && 
b[53038] == 53038 && 
b[53039] == 53039 && 
b[53040] == 53040 && 
b[53041] == 53041 && 
b[53042] == 53042 && 
b[53043] == 53043 && 
b[53044] == 53044 && 
b[53045] == 53045 && 
b[53046] == 53046 && 
b[53047] == 53047 && 
b[53048] == 53048 && 
b[53049] == 53049 && 
b[53050] == 53050 && 
b[53051] == 53051 && 
b[53052] == 53052 && 
b[53053] == 53053 && 
b[53054] == 53054 && 
b[53055] == 53055 && 
b[53056] == 53056 && 
b[53057] == 53057 && 
b[53058] == 53058 && 
b[53059] == 53059 && 
b[53060] == 53060 && 
b[53061] == 53061 && 
b[53062] == 53062 && 
b[53063] == 53063 && 
b[53064] == 53064 && 
b[53065] == 53065 && 
b[53066] == 53066 && 
b[53067] == 53067 && 
b[53068] == 53068 && 
b[53069] == 53069 && 
b[53070] == 53070 && 
b[53071] == 53071 && 
b[53072] == 53072 && 
b[53073] == 53073 && 
b[53074] == 53074 && 
b[53075] == 53075 && 
b[53076] == 53076 && 
b[53077] == 53077 && 
b[53078] == 53078 && 
b[53079] == 53079 && 
b[53080] == 53080 && 
b[53081] == 53081 && 
b[53082] == 53082 && 
b[53083] == 53083 && 
b[53084] == 53084 && 
b[53085] == 53085 && 
b[53086] == 53086 && 
b[53087] == 53087 && 
b[53088] == 53088 && 
b[53089] == 53089 && 
b[53090] == 53090 && 
b[53091] == 53091 && 
b[53092] == 53092 && 
b[53093] == 53093 && 
b[53094] == 53094 && 
b[53095] == 53095 && 
b[53096] == 53096 && 
b[53097] == 53097 && 
b[53098] == 53098 && 
b[53099] == 53099 && 
b[53100] == 53100 && 
b[53101] == 53101 && 
b[53102] == 53102 && 
b[53103] == 53103 && 
b[53104] == 53104 && 
b[53105] == 53105 && 
b[53106] == 53106 && 
b[53107] == 53107 && 
b[53108] == 53108 && 
b[53109] == 53109 && 
b[53110] == 53110 && 
b[53111] == 53111 && 
b[53112] == 53112 && 
b[53113] == 53113 && 
b[53114] == 53114 && 
b[53115] == 53115 && 
b[53116] == 53116 && 
b[53117] == 53117 && 
b[53118] == 53118 && 
b[53119] == 53119 && 
b[53120] == 53120 && 
b[53121] == 53121 && 
b[53122] == 53122 && 
b[53123] == 53123 && 
b[53124] == 53124 && 
b[53125] == 53125 && 
b[53126] == 53126 && 
b[53127] == 53127 && 
b[53128] == 53128 && 
b[53129] == 53129 && 
b[53130] == 53130 && 
b[53131] == 53131 && 
b[53132] == 53132 && 
b[53133] == 53133 && 
b[53134] == 53134 && 
b[53135] == 53135 && 
b[53136] == 53136 && 
b[53137] == 53137 && 
b[53138] == 53138 && 
b[53139] == 53139 && 
b[53140] == 53140 && 
b[53141] == 53141 && 
b[53142] == 53142 && 
b[53143] == 53143 && 
b[53144] == 53144 && 
b[53145] == 53145 && 
b[53146] == 53146 && 
b[53147] == 53147 && 
b[53148] == 53148 && 
b[53149] == 53149 && 
b[53150] == 53150 && 
b[53151] == 53151 && 
b[53152] == 53152 && 
b[53153] == 53153 && 
b[53154] == 53154 && 
b[53155] == 53155 && 
b[53156] == 53156 && 
b[53157] == 53157 && 
b[53158] == 53158 && 
b[53159] == 53159 && 
b[53160] == 53160 && 
b[53161] == 53161 && 
b[53162] == 53162 && 
b[53163] == 53163 && 
b[53164] == 53164 && 
b[53165] == 53165 && 
b[53166] == 53166 && 
b[53167] == 53167 && 
b[53168] == 53168 && 
b[53169] == 53169 && 
b[53170] == 53170 && 
b[53171] == 53171 && 
b[53172] == 53172 && 
b[53173] == 53173 && 
b[53174] == 53174 && 
b[53175] == 53175 && 
b[53176] == 53176 && 
b[53177] == 53177 && 
b[53178] == 53178 && 
b[53179] == 53179 && 
b[53180] == 53180 && 
b[53181] == 53181 && 
b[53182] == 53182 && 
b[53183] == 53183 && 
b[53184] == 53184 && 
b[53185] == 53185 && 
b[53186] == 53186 && 
b[53187] == 53187 && 
b[53188] == 53188 && 
b[53189] == 53189 && 
b[53190] == 53190 && 
b[53191] == 53191 && 
b[53192] == 53192 && 
b[53193] == 53193 && 
b[53194] == 53194 && 
b[53195] == 53195 && 
b[53196] == 53196 && 
b[53197] == 53197 && 
b[53198] == 53198 && 
b[53199] == 53199 && 
b[53200] == 53200 && 
b[53201] == 53201 && 
b[53202] == 53202 && 
b[53203] == 53203 && 
b[53204] == 53204 && 
b[53205] == 53205 && 
b[53206] == 53206 && 
b[53207] == 53207 && 
b[53208] == 53208 && 
b[53209] == 53209 && 
b[53210] == 53210 && 
b[53211] == 53211 && 
b[53212] == 53212 && 
b[53213] == 53213 && 
b[53214] == 53214 && 
b[53215] == 53215 && 
b[53216] == 53216 && 
b[53217] == 53217 && 
b[53218] == 53218 && 
b[53219] == 53219 && 
b[53220] == 53220 && 
b[53221] == 53221 && 
b[53222] == 53222 && 
b[53223] == 53223 && 
b[53224] == 53224 && 
b[53225] == 53225 && 
b[53226] == 53226 && 
b[53227] == 53227 && 
b[53228] == 53228 && 
b[53229] == 53229 && 
b[53230] == 53230 && 
b[53231] == 53231 && 
b[53232] == 53232 && 
b[53233] == 53233 && 
b[53234] == 53234 && 
b[53235] == 53235 && 
b[53236] == 53236 && 
b[53237] == 53237 && 
b[53238] == 53238 && 
b[53239] == 53239 && 
b[53240] == 53240 && 
b[53241] == 53241 && 
b[53242] == 53242 && 
b[53243] == 53243 && 
b[53244] == 53244 && 
b[53245] == 53245 && 
b[53246] == 53246 && 
b[53247] == 53247 && 
b[53248] == 53248 && 
b[53249] == 53249 && 
b[53250] == 53250 && 
b[53251] == 53251 && 
b[53252] == 53252 && 
b[53253] == 53253 && 
b[53254] == 53254 && 
b[53255] == 53255 && 
b[53256] == 53256 && 
b[53257] == 53257 && 
b[53258] == 53258 && 
b[53259] == 53259 && 
b[53260] == 53260 && 
b[53261] == 53261 && 
b[53262] == 53262 && 
b[53263] == 53263 && 
b[53264] == 53264 && 
b[53265] == 53265 && 
b[53266] == 53266 && 
b[53267] == 53267 && 
b[53268] == 53268 && 
b[53269] == 53269 && 
b[53270] == 53270 && 
b[53271] == 53271 && 
b[53272] == 53272 && 
b[53273] == 53273 && 
b[53274] == 53274 && 
b[53275] == 53275 && 
b[53276] == 53276 && 
b[53277] == 53277 && 
b[53278] == 53278 && 
b[53279] == 53279 && 
b[53280] == 53280 && 
b[53281] == 53281 && 
b[53282] == 53282 && 
b[53283] == 53283 && 
b[53284] == 53284 && 
b[53285] == 53285 && 
b[53286] == 53286 && 
b[53287] == 53287 && 
b[53288] == 53288 && 
b[53289] == 53289 && 
b[53290] == 53290 && 
b[53291] == 53291 && 
b[53292] == 53292 && 
b[53293] == 53293 && 
b[53294] == 53294 && 
b[53295] == 53295 && 
b[53296] == 53296 && 
b[53297] == 53297 && 
b[53298] == 53298 && 
b[53299] == 53299 && 
b[53300] == 53300 && 
b[53301] == 53301 && 
b[53302] == 53302 && 
b[53303] == 53303 && 
b[53304] == 53304 && 
b[53305] == 53305 && 
b[53306] == 53306 && 
b[53307] == 53307 && 
b[53308] == 53308 && 
b[53309] == 53309 && 
b[53310] == 53310 && 
b[53311] == 53311 && 
b[53312] == 53312 && 
b[53313] == 53313 && 
b[53314] == 53314 && 
b[53315] == 53315 && 
b[53316] == 53316 && 
b[53317] == 53317 && 
b[53318] == 53318 && 
b[53319] == 53319 && 
b[53320] == 53320 && 
b[53321] == 53321 && 
b[53322] == 53322 && 
b[53323] == 53323 && 
b[53324] == 53324 && 
b[53325] == 53325 && 
b[53326] == 53326 && 
b[53327] == 53327 && 
b[53328] == 53328 && 
b[53329] == 53329 && 
b[53330] == 53330 && 
b[53331] == 53331 && 
b[53332] == 53332 && 
b[53333] == 53333 && 
b[53334] == 53334 && 
b[53335] == 53335 && 
b[53336] == 53336 && 
b[53337] == 53337 && 
b[53338] == 53338 && 
b[53339] == 53339 && 
b[53340] == 53340 && 
b[53341] == 53341 && 
b[53342] == 53342 && 
b[53343] == 53343 && 
b[53344] == 53344 && 
b[53345] == 53345 && 
b[53346] == 53346 && 
b[53347] == 53347 && 
b[53348] == 53348 && 
b[53349] == 53349 && 
b[53350] == 53350 && 
b[53351] == 53351 && 
b[53352] == 53352 && 
b[53353] == 53353 && 
b[53354] == 53354 && 
b[53355] == 53355 && 
b[53356] == 53356 && 
b[53357] == 53357 && 
b[53358] == 53358 && 
b[53359] == 53359 && 
b[53360] == 53360 && 
b[53361] == 53361 && 
b[53362] == 53362 && 
b[53363] == 53363 && 
b[53364] == 53364 && 
b[53365] == 53365 && 
b[53366] == 53366 && 
b[53367] == 53367 && 
b[53368] == 53368 && 
b[53369] == 53369 && 
b[53370] == 53370 && 
b[53371] == 53371 && 
b[53372] == 53372 && 
b[53373] == 53373 && 
b[53374] == 53374 && 
b[53375] == 53375 && 
b[53376] == 53376 && 
b[53377] == 53377 && 
b[53378] == 53378 && 
b[53379] == 53379 && 
b[53380] == 53380 && 
b[53381] == 53381 && 
b[53382] == 53382 && 
b[53383] == 53383 && 
b[53384] == 53384 && 
b[53385] == 53385 && 
b[53386] == 53386 && 
b[53387] == 53387 && 
b[53388] == 53388 && 
b[53389] == 53389 && 
b[53390] == 53390 && 
b[53391] == 53391 && 
b[53392] == 53392 && 
b[53393] == 53393 && 
b[53394] == 53394 && 
b[53395] == 53395 && 
b[53396] == 53396 && 
b[53397] == 53397 && 
b[53398] == 53398 && 
b[53399] == 53399 && 
b[53400] == 53400 && 
b[53401] == 53401 && 
b[53402] == 53402 && 
b[53403] == 53403 && 
b[53404] == 53404 && 
b[53405] == 53405 && 
b[53406] == 53406 && 
b[53407] == 53407 && 
b[53408] == 53408 && 
b[53409] == 53409 && 
b[53410] == 53410 && 
b[53411] == 53411 && 
b[53412] == 53412 && 
b[53413] == 53413 && 
b[53414] == 53414 && 
b[53415] == 53415 && 
b[53416] == 53416 && 
b[53417] == 53417 && 
b[53418] == 53418 && 
b[53419] == 53419 && 
b[53420] == 53420 && 
b[53421] == 53421 && 
b[53422] == 53422 && 
b[53423] == 53423 && 
b[53424] == 53424 && 
b[53425] == 53425 && 
b[53426] == 53426 && 
b[53427] == 53427 && 
b[53428] == 53428 && 
b[53429] == 53429 && 
b[53430] == 53430 && 
b[53431] == 53431 && 
b[53432] == 53432 && 
b[53433] == 53433 && 
b[53434] == 53434 && 
b[53435] == 53435 && 
b[53436] == 53436 && 
b[53437] == 53437 && 
b[53438] == 53438 && 
b[53439] == 53439 && 
b[53440] == 53440 && 
b[53441] == 53441 && 
b[53442] == 53442 && 
b[53443] == 53443 && 
b[53444] == 53444 && 
b[53445] == 53445 && 
b[53446] == 53446 && 
b[53447] == 53447 && 
b[53448] == 53448 && 
b[53449] == 53449 && 
b[53450] == 53450 && 
b[53451] == 53451 && 
b[53452] == 53452 && 
b[53453] == 53453 && 
b[53454] == 53454 && 
b[53455] == 53455 && 
b[53456] == 53456 && 
b[53457] == 53457 && 
b[53458] == 53458 && 
b[53459] == 53459 && 
b[53460] == 53460 && 
b[53461] == 53461 && 
b[53462] == 53462 && 
b[53463] == 53463 && 
b[53464] == 53464 && 
b[53465] == 53465 && 
b[53466] == 53466 && 
b[53467] == 53467 && 
b[53468] == 53468 && 
b[53469] == 53469 && 
b[53470] == 53470 && 
b[53471] == 53471 && 
b[53472] == 53472 && 
b[53473] == 53473 && 
b[53474] == 53474 && 
b[53475] == 53475 && 
b[53476] == 53476 && 
b[53477] == 53477 && 
b[53478] == 53478 && 
b[53479] == 53479 && 
b[53480] == 53480 && 
b[53481] == 53481 && 
b[53482] == 53482 && 
b[53483] == 53483 && 
b[53484] == 53484 && 
b[53485] == 53485 && 
b[53486] == 53486 && 
b[53487] == 53487 && 
b[53488] == 53488 && 
b[53489] == 53489 && 
b[53490] == 53490 && 
b[53491] == 53491 && 
b[53492] == 53492 && 
b[53493] == 53493 && 
b[53494] == 53494 && 
b[53495] == 53495 && 
b[53496] == 53496 && 
b[53497] == 53497 && 
b[53498] == 53498 && 
b[53499] == 53499 && 
b[53500] == 53500 && 
b[53501] == 53501 && 
b[53502] == 53502 && 
b[53503] == 53503 && 
b[53504] == 53504 && 
b[53505] == 53505 && 
b[53506] == 53506 && 
b[53507] == 53507 && 
b[53508] == 53508 && 
b[53509] == 53509 && 
b[53510] == 53510 && 
b[53511] == 53511 && 
b[53512] == 53512 && 
b[53513] == 53513 && 
b[53514] == 53514 && 
b[53515] == 53515 && 
b[53516] == 53516 && 
b[53517] == 53517 && 
b[53518] == 53518 && 
b[53519] == 53519 && 
b[53520] == 53520 && 
b[53521] == 53521 && 
b[53522] == 53522 && 
b[53523] == 53523 && 
b[53524] == 53524 && 
b[53525] == 53525 && 
b[53526] == 53526 && 
b[53527] == 53527 && 
b[53528] == 53528 && 
b[53529] == 53529 && 
b[53530] == 53530 && 
b[53531] == 53531 && 
b[53532] == 53532 && 
b[53533] == 53533 && 
b[53534] == 53534 && 
b[53535] == 53535 && 
b[53536] == 53536 && 
b[53537] == 53537 && 
b[53538] == 53538 && 
b[53539] == 53539 && 
b[53540] == 53540 && 
b[53541] == 53541 && 
b[53542] == 53542 && 
b[53543] == 53543 && 
b[53544] == 53544 && 
b[53545] == 53545 && 
b[53546] == 53546 && 
b[53547] == 53547 && 
b[53548] == 53548 && 
b[53549] == 53549 && 
b[53550] == 53550 && 
b[53551] == 53551 && 
b[53552] == 53552 && 
b[53553] == 53553 && 
b[53554] == 53554 && 
b[53555] == 53555 && 
b[53556] == 53556 && 
b[53557] == 53557 && 
b[53558] == 53558 && 
b[53559] == 53559 && 
b[53560] == 53560 && 
b[53561] == 53561 && 
b[53562] == 53562 && 
b[53563] == 53563 && 
b[53564] == 53564 && 
b[53565] == 53565 && 
b[53566] == 53566 && 
b[53567] == 53567 && 
b[53568] == 53568 && 
b[53569] == 53569 && 
b[53570] == 53570 && 
b[53571] == 53571 && 
b[53572] == 53572 && 
b[53573] == 53573 && 
b[53574] == 53574 && 
b[53575] == 53575 && 
b[53576] == 53576 && 
b[53577] == 53577 && 
b[53578] == 53578 && 
b[53579] == 53579 && 
b[53580] == 53580 && 
b[53581] == 53581 && 
b[53582] == 53582 && 
b[53583] == 53583 && 
b[53584] == 53584 && 
b[53585] == 53585 && 
b[53586] == 53586 && 
b[53587] == 53587 && 
b[53588] == 53588 && 
b[53589] == 53589 && 
b[53590] == 53590 && 
b[53591] == 53591 && 
b[53592] == 53592 && 
b[53593] == 53593 && 
b[53594] == 53594 && 
b[53595] == 53595 && 
b[53596] == 53596 && 
b[53597] == 53597 && 
b[53598] == 53598 && 
b[53599] == 53599 && 
b[53600] == 53600 && 
b[53601] == 53601 && 
b[53602] == 53602 && 
b[53603] == 53603 && 
b[53604] == 53604 && 
b[53605] == 53605 && 
b[53606] == 53606 && 
b[53607] == 53607 && 
b[53608] == 53608 && 
b[53609] == 53609 && 
b[53610] == 53610 && 
b[53611] == 53611 && 
b[53612] == 53612 && 
b[53613] == 53613 && 
b[53614] == 53614 && 
b[53615] == 53615 && 
b[53616] == 53616 && 
b[53617] == 53617 && 
b[53618] == 53618 && 
b[53619] == 53619 && 
b[53620] == 53620 && 
b[53621] == 53621 && 
b[53622] == 53622 && 
b[53623] == 53623 && 
b[53624] == 53624 && 
b[53625] == 53625 && 
b[53626] == 53626 && 
b[53627] == 53627 && 
b[53628] == 53628 && 
b[53629] == 53629 && 
b[53630] == 53630 && 
b[53631] == 53631 && 
b[53632] == 53632 && 
b[53633] == 53633 && 
b[53634] == 53634 && 
b[53635] == 53635 && 
b[53636] == 53636 && 
b[53637] == 53637 && 
b[53638] == 53638 && 
b[53639] == 53639 && 
b[53640] == 53640 && 
b[53641] == 53641 && 
b[53642] == 53642 && 
b[53643] == 53643 && 
b[53644] == 53644 && 
b[53645] == 53645 && 
b[53646] == 53646 && 
b[53647] == 53647 && 
b[53648] == 53648 && 
b[53649] == 53649 && 
b[53650] == 53650 && 
b[53651] == 53651 && 
b[53652] == 53652 && 
b[53653] == 53653 && 
b[53654] == 53654 && 
b[53655] == 53655 && 
b[53656] == 53656 && 
b[53657] == 53657 && 
b[53658] == 53658 && 
b[53659] == 53659 && 
b[53660] == 53660 && 
b[53661] == 53661 && 
b[53662] == 53662 && 
b[53663] == 53663 && 
b[53664] == 53664 && 
b[53665] == 53665 && 
b[53666] == 53666 && 
b[53667] == 53667 && 
b[53668] == 53668 && 
b[53669] == 53669 && 
b[53670] == 53670 && 
b[53671] == 53671 && 
b[53672] == 53672 && 
b[53673] == 53673 && 
b[53674] == 53674 && 
b[53675] == 53675 && 
b[53676] == 53676 && 
b[53677] == 53677 && 
b[53678] == 53678 && 
b[53679] == 53679 && 
b[53680] == 53680 && 
b[53681] == 53681 && 
b[53682] == 53682 && 
b[53683] == 53683 && 
b[53684] == 53684 && 
b[53685] == 53685 && 
b[53686] == 53686 && 
b[53687] == 53687 && 
b[53688] == 53688 && 
b[53689] == 53689 && 
b[53690] == 53690 && 
b[53691] == 53691 && 
b[53692] == 53692 && 
b[53693] == 53693 && 
b[53694] == 53694 && 
b[53695] == 53695 && 
b[53696] == 53696 && 
b[53697] == 53697 && 
b[53698] == 53698 && 
b[53699] == 53699 && 
b[53700] == 53700 && 
b[53701] == 53701 && 
b[53702] == 53702 && 
b[53703] == 53703 && 
b[53704] == 53704 && 
b[53705] == 53705 && 
b[53706] == 53706 && 
b[53707] == 53707 && 
b[53708] == 53708 && 
b[53709] == 53709 && 
b[53710] == 53710 && 
b[53711] == 53711 && 
b[53712] == 53712 && 
b[53713] == 53713 && 
b[53714] == 53714 && 
b[53715] == 53715 && 
b[53716] == 53716 && 
b[53717] == 53717 && 
b[53718] == 53718 && 
b[53719] == 53719 && 
b[53720] == 53720 && 
b[53721] == 53721 && 
b[53722] == 53722 && 
b[53723] == 53723 && 
b[53724] == 53724 && 
b[53725] == 53725 && 
b[53726] == 53726 && 
b[53727] == 53727 && 
b[53728] == 53728 && 
b[53729] == 53729 && 
b[53730] == 53730 && 
b[53731] == 53731 && 
b[53732] == 53732 && 
b[53733] == 53733 && 
b[53734] == 53734 && 
b[53735] == 53735 && 
b[53736] == 53736 && 
b[53737] == 53737 && 
b[53738] == 53738 && 
b[53739] == 53739 && 
b[53740] == 53740 && 
b[53741] == 53741 && 
b[53742] == 53742 && 
b[53743] == 53743 && 
b[53744] == 53744 && 
b[53745] == 53745 && 
b[53746] == 53746 && 
b[53747] == 53747 && 
b[53748] == 53748 && 
b[53749] == 53749 && 
b[53750] == 53750 && 
b[53751] == 53751 && 
b[53752] == 53752 && 
b[53753] == 53753 && 
b[53754] == 53754 && 
b[53755] == 53755 && 
b[53756] == 53756 && 
b[53757] == 53757 && 
b[53758] == 53758 && 
b[53759] == 53759 && 
b[53760] == 53760 && 
b[53761] == 53761 && 
b[53762] == 53762 && 
b[53763] == 53763 && 
b[53764] == 53764 && 
b[53765] == 53765 && 
b[53766] == 53766 && 
b[53767] == 53767 && 
b[53768] == 53768 && 
b[53769] == 53769 && 
b[53770] == 53770 && 
b[53771] == 53771 && 
b[53772] == 53772 && 
b[53773] == 53773 && 
b[53774] == 53774 && 
b[53775] == 53775 && 
b[53776] == 53776 && 
b[53777] == 53777 && 
b[53778] == 53778 && 
b[53779] == 53779 && 
b[53780] == 53780 && 
b[53781] == 53781 && 
b[53782] == 53782 && 
b[53783] == 53783 && 
b[53784] == 53784 && 
b[53785] == 53785 && 
b[53786] == 53786 && 
b[53787] == 53787 && 
b[53788] == 53788 && 
b[53789] == 53789 && 
b[53790] == 53790 && 
b[53791] == 53791 && 
b[53792] == 53792 && 
b[53793] == 53793 && 
b[53794] == 53794 && 
b[53795] == 53795 && 
b[53796] == 53796 && 
b[53797] == 53797 && 
b[53798] == 53798 && 
b[53799] == 53799 && 
b[53800] == 53800 && 
b[53801] == 53801 && 
b[53802] == 53802 && 
b[53803] == 53803 && 
b[53804] == 53804 && 
b[53805] == 53805 && 
b[53806] == 53806 && 
b[53807] == 53807 && 
b[53808] == 53808 && 
b[53809] == 53809 && 
b[53810] == 53810 && 
b[53811] == 53811 && 
b[53812] == 53812 && 
b[53813] == 53813 && 
b[53814] == 53814 && 
b[53815] == 53815 && 
b[53816] == 53816 && 
b[53817] == 53817 && 
b[53818] == 53818 && 
b[53819] == 53819 && 
b[53820] == 53820 && 
b[53821] == 53821 && 
b[53822] == 53822 && 
b[53823] == 53823 && 
b[53824] == 53824 && 
b[53825] == 53825 && 
b[53826] == 53826 && 
b[53827] == 53827 && 
b[53828] == 53828 && 
b[53829] == 53829 && 
b[53830] == 53830 && 
b[53831] == 53831 && 
b[53832] == 53832 && 
b[53833] == 53833 && 
b[53834] == 53834 && 
b[53835] == 53835 && 
b[53836] == 53836 && 
b[53837] == 53837 && 
b[53838] == 53838 && 
b[53839] == 53839 && 
b[53840] == 53840 && 
b[53841] == 53841 && 
b[53842] == 53842 && 
b[53843] == 53843 && 
b[53844] == 53844 && 
b[53845] == 53845 && 
b[53846] == 53846 && 
b[53847] == 53847 && 
b[53848] == 53848 && 
b[53849] == 53849 && 
b[53850] == 53850 && 
b[53851] == 53851 && 
b[53852] == 53852 && 
b[53853] == 53853 && 
b[53854] == 53854 && 
b[53855] == 53855 && 
b[53856] == 53856 && 
b[53857] == 53857 && 
b[53858] == 53858 && 
b[53859] == 53859 && 
b[53860] == 53860 && 
b[53861] == 53861 && 
b[53862] == 53862 && 
b[53863] == 53863 && 
b[53864] == 53864 && 
b[53865] == 53865 && 
b[53866] == 53866 && 
b[53867] == 53867 && 
b[53868] == 53868 && 
b[53869] == 53869 && 
b[53870] == 53870 && 
b[53871] == 53871 && 
b[53872] == 53872 && 
b[53873] == 53873 && 
b[53874] == 53874 && 
b[53875] == 53875 && 
b[53876] == 53876 && 
b[53877] == 53877 && 
b[53878] == 53878 && 
b[53879] == 53879 && 
b[53880] == 53880 && 
b[53881] == 53881 && 
b[53882] == 53882 && 
b[53883] == 53883 && 
b[53884] == 53884 && 
b[53885] == 53885 && 
b[53886] == 53886 && 
b[53887] == 53887 && 
b[53888] == 53888 && 
b[53889] == 53889 && 
b[53890] == 53890 && 
b[53891] == 53891 && 
b[53892] == 53892 && 
b[53893] == 53893 && 
b[53894] == 53894 && 
b[53895] == 53895 && 
b[53896] == 53896 && 
b[53897] == 53897 && 
b[53898] == 53898 && 
b[53899] == 53899 && 
b[53900] == 53900 && 
b[53901] == 53901 && 
b[53902] == 53902 && 
b[53903] == 53903 && 
b[53904] == 53904 && 
b[53905] == 53905 && 
b[53906] == 53906 && 
b[53907] == 53907 && 
b[53908] == 53908 && 
b[53909] == 53909 && 
b[53910] == 53910 && 
b[53911] == 53911 && 
b[53912] == 53912 && 
b[53913] == 53913 && 
b[53914] == 53914 && 
b[53915] == 53915 && 
b[53916] == 53916 && 
b[53917] == 53917 && 
b[53918] == 53918 && 
b[53919] == 53919 && 
b[53920] == 53920 && 
b[53921] == 53921 && 
b[53922] == 53922 && 
b[53923] == 53923 && 
b[53924] == 53924 && 
b[53925] == 53925 && 
b[53926] == 53926 && 
b[53927] == 53927 && 
b[53928] == 53928 && 
b[53929] == 53929 && 
b[53930] == 53930 && 
b[53931] == 53931 && 
b[53932] == 53932 && 
b[53933] == 53933 && 
b[53934] == 53934 && 
b[53935] == 53935 && 
b[53936] == 53936 && 
b[53937] == 53937 && 
b[53938] == 53938 && 
b[53939] == 53939 && 
b[53940] == 53940 && 
b[53941] == 53941 && 
b[53942] == 53942 && 
b[53943] == 53943 && 
b[53944] == 53944 && 
b[53945] == 53945 && 
b[53946] == 53946 && 
b[53947] == 53947 && 
b[53948] == 53948 && 
b[53949] == 53949 && 
b[53950] == 53950 && 
b[53951] == 53951 && 
b[53952] == 53952 && 
b[53953] == 53953 && 
b[53954] == 53954 && 
b[53955] == 53955 && 
b[53956] == 53956 && 
b[53957] == 53957 && 
b[53958] == 53958 && 
b[53959] == 53959 && 
b[53960] == 53960 && 
b[53961] == 53961 && 
b[53962] == 53962 && 
b[53963] == 53963 && 
b[53964] == 53964 && 
b[53965] == 53965 && 
b[53966] == 53966 && 
b[53967] == 53967 && 
b[53968] == 53968 && 
b[53969] == 53969 && 
b[53970] == 53970 && 
b[53971] == 53971 && 
b[53972] == 53972 && 
b[53973] == 53973 && 
b[53974] == 53974 && 
b[53975] == 53975 && 
b[53976] == 53976 && 
b[53977] == 53977 && 
b[53978] == 53978 && 
b[53979] == 53979 && 
b[53980] == 53980 && 
b[53981] == 53981 && 
b[53982] == 53982 && 
b[53983] == 53983 && 
b[53984] == 53984 && 
b[53985] == 53985 && 
b[53986] == 53986 && 
b[53987] == 53987 && 
b[53988] == 53988 && 
b[53989] == 53989 && 
b[53990] == 53990 && 
b[53991] == 53991 && 
b[53992] == 53992 && 
b[53993] == 53993 && 
b[53994] == 53994 && 
b[53995] == 53995 && 
b[53996] == 53996 && 
b[53997] == 53997 && 
b[53998] == 53998 && 
b[53999] == 53999 && 
b[54000] == 54000 && 
b[54001] == 54001 && 
b[54002] == 54002 && 
b[54003] == 54003 && 
b[54004] == 54004 && 
b[54005] == 54005 && 
b[54006] == 54006 && 
b[54007] == 54007 && 
b[54008] == 54008 && 
b[54009] == 54009 && 
b[54010] == 54010 && 
b[54011] == 54011 && 
b[54012] == 54012 && 
b[54013] == 54013 && 
b[54014] == 54014 && 
b[54015] == 54015 && 
b[54016] == 54016 && 
b[54017] == 54017 && 
b[54018] == 54018 && 
b[54019] == 54019 && 
b[54020] == 54020 && 
b[54021] == 54021 && 
b[54022] == 54022 && 
b[54023] == 54023 && 
b[54024] == 54024 && 
b[54025] == 54025 && 
b[54026] == 54026 && 
b[54027] == 54027 && 
b[54028] == 54028 && 
b[54029] == 54029 && 
b[54030] == 54030 && 
b[54031] == 54031 && 
b[54032] == 54032 && 
b[54033] == 54033 && 
b[54034] == 54034 && 
b[54035] == 54035 && 
b[54036] == 54036 && 
b[54037] == 54037 && 
b[54038] == 54038 && 
b[54039] == 54039 && 
b[54040] == 54040 && 
b[54041] == 54041 && 
b[54042] == 54042 && 
b[54043] == 54043 && 
b[54044] == 54044 && 
b[54045] == 54045 && 
b[54046] == 54046 && 
b[54047] == 54047 && 
b[54048] == 54048 && 
b[54049] == 54049 && 
b[54050] == 54050 && 
b[54051] == 54051 && 
b[54052] == 54052 && 
b[54053] == 54053 && 
b[54054] == 54054 && 
b[54055] == 54055 && 
b[54056] == 54056 && 
b[54057] == 54057 && 
b[54058] == 54058 && 
b[54059] == 54059 && 
b[54060] == 54060 && 
b[54061] == 54061 && 
b[54062] == 54062 && 
b[54063] == 54063 && 
b[54064] == 54064 && 
b[54065] == 54065 && 
b[54066] == 54066 && 
b[54067] == 54067 && 
b[54068] == 54068 && 
b[54069] == 54069 && 
b[54070] == 54070 && 
b[54071] == 54071 && 
b[54072] == 54072 && 
b[54073] == 54073 && 
b[54074] == 54074 && 
b[54075] == 54075 && 
b[54076] == 54076 && 
b[54077] == 54077 && 
b[54078] == 54078 && 
b[54079] == 54079 && 
b[54080] == 54080 && 
b[54081] == 54081 && 
b[54082] == 54082 && 
b[54083] == 54083 && 
b[54084] == 54084 && 
b[54085] == 54085 && 
b[54086] == 54086 && 
b[54087] == 54087 && 
b[54088] == 54088 && 
b[54089] == 54089 && 
b[54090] == 54090 && 
b[54091] == 54091 && 
b[54092] == 54092 && 
b[54093] == 54093 && 
b[54094] == 54094 && 
b[54095] == 54095 && 
b[54096] == 54096 && 
b[54097] == 54097 && 
b[54098] == 54098 && 
b[54099] == 54099 && 
b[54100] == 54100 && 
b[54101] == 54101 && 
b[54102] == 54102 && 
b[54103] == 54103 && 
b[54104] == 54104 && 
b[54105] == 54105 && 
b[54106] == 54106 && 
b[54107] == 54107 && 
b[54108] == 54108 && 
b[54109] == 54109 && 
b[54110] == 54110 && 
b[54111] == 54111 && 
b[54112] == 54112 && 
b[54113] == 54113 && 
b[54114] == 54114 && 
b[54115] == 54115 && 
b[54116] == 54116 && 
b[54117] == 54117 && 
b[54118] == 54118 && 
b[54119] == 54119 && 
b[54120] == 54120 && 
b[54121] == 54121 && 
b[54122] == 54122 && 
b[54123] == 54123 && 
b[54124] == 54124 && 
b[54125] == 54125 && 
b[54126] == 54126 && 
b[54127] == 54127 && 
b[54128] == 54128 && 
b[54129] == 54129 && 
b[54130] == 54130 && 
b[54131] == 54131 && 
b[54132] == 54132 && 
b[54133] == 54133 && 
b[54134] == 54134 && 
b[54135] == 54135 && 
b[54136] == 54136 && 
b[54137] == 54137 && 
b[54138] == 54138 && 
b[54139] == 54139 && 
b[54140] == 54140 && 
b[54141] == 54141 && 
b[54142] == 54142 && 
b[54143] == 54143 && 
b[54144] == 54144 && 
b[54145] == 54145 && 
b[54146] == 54146 && 
b[54147] == 54147 && 
b[54148] == 54148 && 
b[54149] == 54149 && 
b[54150] == 54150 && 
b[54151] == 54151 && 
b[54152] == 54152 && 
b[54153] == 54153 && 
b[54154] == 54154 && 
b[54155] == 54155 && 
b[54156] == 54156 && 
b[54157] == 54157 && 
b[54158] == 54158 && 
b[54159] == 54159 && 
b[54160] == 54160 && 
b[54161] == 54161 && 
b[54162] == 54162 && 
b[54163] == 54163 && 
b[54164] == 54164 && 
b[54165] == 54165 && 
b[54166] == 54166 && 
b[54167] == 54167 && 
b[54168] == 54168 && 
b[54169] == 54169 && 
b[54170] == 54170 && 
b[54171] == 54171 && 
b[54172] == 54172 && 
b[54173] == 54173 && 
b[54174] == 54174 && 
b[54175] == 54175 && 
b[54176] == 54176 && 
b[54177] == 54177 && 
b[54178] == 54178 && 
b[54179] == 54179 && 
b[54180] == 54180 && 
b[54181] == 54181 && 
b[54182] == 54182 && 
b[54183] == 54183 && 
b[54184] == 54184 && 
b[54185] == 54185 && 
b[54186] == 54186 && 
b[54187] == 54187 && 
b[54188] == 54188 && 
b[54189] == 54189 && 
b[54190] == 54190 && 
b[54191] == 54191 && 
b[54192] == 54192 && 
b[54193] == 54193 && 
b[54194] == 54194 && 
b[54195] == 54195 && 
b[54196] == 54196 && 
b[54197] == 54197 && 
b[54198] == 54198 && 
b[54199] == 54199 && 
b[54200] == 54200 && 
b[54201] == 54201 && 
b[54202] == 54202 && 
b[54203] == 54203 && 
b[54204] == 54204 && 
b[54205] == 54205 && 
b[54206] == 54206 && 
b[54207] == 54207 && 
b[54208] == 54208 && 
b[54209] == 54209 && 
b[54210] == 54210 && 
b[54211] == 54211 && 
b[54212] == 54212 && 
b[54213] == 54213 && 
b[54214] == 54214 && 
b[54215] == 54215 && 
b[54216] == 54216 && 
b[54217] == 54217 && 
b[54218] == 54218 && 
b[54219] == 54219 && 
b[54220] == 54220 && 
b[54221] == 54221 && 
b[54222] == 54222 && 
b[54223] == 54223 && 
b[54224] == 54224 && 
b[54225] == 54225 && 
b[54226] == 54226 && 
b[54227] == 54227 && 
b[54228] == 54228 && 
b[54229] == 54229 && 
b[54230] == 54230 && 
b[54231] == 54231 && 
b[54232] == 54232 && 
b[54233] == 54233 && 
b[54234] == 54234 && 
b[54235] == 54235 && 
b[54236] == 54236 && 
b[54237] == 54237 && 
b[54238] == 54238 && 
b[54239] == 54239 && 
b[54240] == 54240 && 
b[54241] == 54241 && 
b[54242] == 54242 && 
b[54243] == 54243 && 
b[54244] == 54244 && 
b[54245] == 54245 && 
b[54246] == 54246 && 
b[54247] == 54247 && 
b[54248] == 54248 && 
b[54249] == 54249 && 
b[54250] == 54250 && 
b[54251] == 54251 && 
b[54252] == 54252 && 
b[54253] == 54253 && 
b[54254] == 54254 && 
b[54255] == 54255 && 
b[54256] == 54256 && 
b[54257] == 54257 && 
b[54258] == 54258 && 
b[54259] == 54259 && 
b[54260] == 54260 && 
b[54261] == 54261 && 
b[54262] == 54262 && 
b[54263] == 54263 && 
b[54264] == 54264 && 
b[54265] == 54265 && 
b[54266] == 54266 && 
b[54267] == 54267 && 
b[54268] == 54268 && 
b[54269] == 54269 && 
b[54270] == 54270 && 
b[54271] == 54271 && 
b[54272] == 54272 && 
b[54273] == 54273 && 
b[54274] == 54274 && 
b[54275] == 54275 && 
b[54276] == 54276 && 
b[54277] == 54277 && 
b[54278] == 54278 && 
b[54279] == 54279 && 
b[54280] == 54280 && 
b[54281] == 54281 && 
b[54282] == 54282 && 
b[54283] == 54283 && 
b[54284] == 54284 && 
b[54285] == 54285 && 
b[54286] == 54286 && 
b[54287] == 54287 && 
b[54288] == 54288 && 
b[54289] == 54289 && 
b[54290] == 54290 && 
b[54291] == 54291 && 
b[54292] == 54292 && 
b[54293] == 54293 && 
b[54294] == 54294 && 
b[54295] == 54295 && 
b[54296] == 54296 && 
b[54297] == 54297 && 
b[54298] == 54298 && 
b[54299] == 54299 && 
b[54300] == 54300 && 
b[54301] == 54301 && 
b[54302] == 54302 && 
b[54303] == 54303 && 
b[54304] == 54304 && 
b[54305] == 54305 && 
b[54306] == 54306 && 
b[54307] == 54307 && 
b[54308] == 54308 && 
b[54309] == 54309 && 
b[54310] == 54310 && 
b[54311] == 54311 && 
b[54312] == 54312 && 
b[54313] == 54313 && 
b[54314] == 54314 && 
b[54315] == 54315 && 
b[54316] == 54316 && 
b[54317] == 54317 && 
b[54318] == 54318 && 
b[54319] == 54319 && 
b[54320] == 54320 && 
b[54321] == 54321 && 
b[54322] == 54322 && 
b[54323] == 54323 && 
b[54324] == 54324 && 
b[54325] == 54325 && 
b[54326] == 54326 && 
b[54327] == 54327 && 
b[54328] == 54328 && 
b[54329] == 54329 && 
b[54330] == 54330 && 
b[54331] == 54331 && 
b[54332] == 54332 && 
b[54333] == 54333 && 
b[54334] == 54334 && 
b[54335] == 54335 && 
b[54336] == 54336 && 
b[54337] == 54337 && 
b[54338] == 54338 && 
b[54339] == 54339 && 
b[54340] == 54340 && 
b[54341] == 54341 && 
b[54342] == 54342 && 
b[54343] == 54343 && 
b[54344] == 54344 && 
b[54345] == 54345 && 
b[54346] == 54346 && 
b[54347] == 54347 && 
b[54348] == 54348 && 
b[54349] == 54349 && 
b[54350] == 54350 && 
b[54351] == 54351 && 
b[54352] == 54352 && 
b[54353] == 54353 && 
b[54354] == 54354 && 
b[54355] == 54355 && 
b[54356] == 54356 && 
b[54357] == 54357 && 
b[54358] == 54358 && 
b[54359] == 54359 && 
b[54360] == 54360 && 
b[54361] == 54361 && 
b[54362] == 54362 && 
b[54363] == 54363 && 
b[54364] == 54364 && 
b[54365] == 54365 && 
b[54366] == 54366 && 
b[54367] == 54367 && 
b[54368] == 54368 && 
b[54369] == 54369 && 
b[54370] == 54370 && 
b[54371] == 54371 && 
b[54372] == 54372 && 
b[54373] == 54373 && 
b[54374] == 54374 && 
b[54375] == 54375 && 
b[54376] == 54376 && 
b[54377] == 54377 && 
b[54378] == 54378 && 
b[54379] == 54379 && 
b[54380] == 54380 && 
b[54381] == 54381 && 
b[54382] == 54382 && 
b[54383] == 54383 && 
b[54384] == 54384 && 
b[54385] == 54385 && 
b[54386] == 54386 && 
b[54387] == 54387 && 
b[54388] == 54388 && 
b[54389] == 54389 && 
b[54390] == 54390 && 
b[54391] == 54391 && 
b[54392] == 54392 && 
b[54393] == 54393 && 
b[54394] == 54394 && 
b[54395] == 54395 && 
b[54396] == 54396 && 
b[54397] == 54397 && 
b[54398] == 54398 && 
b[54399] == 54399 && 
b[54400] == 54400 && 
b[54401] == 54401 && 
b[54402] == 54402 && 
b[54403] == 54403 && 
b[54404] == 54404 && 
b[54405] == 54405 && 
b[54406] == 54406 && 
b[54407] == 54407 && 
b[54408] == 54408 && 
b[54409] == 54409 && 
b[54410] == 54410 && 
b[54411] == 54411 && 
b[54412] == 54412 && 
b[54413] == 54413 && 
b[54414] == 54414 && 
b[54415] == 54415 && 
b[54416] == 54416 && 
b[54417] == 54417 && 
b[54418] == 54418 && 
b[54419] == 54419 && 
b[54420] == 54420 && 
b[54421] == 54421 && 
b[54422] == 54422 && 
b[54423] == 54423 && 
b[54424] == 54424 && 
b[54425] == 54425 && 
b[54426] == 54426 && 
b[54427] == 54427 && 
b[54428] == 54428 && 
b[54429] == 54429 && 
b[54430] == 54430 && 
b[54431] == 54431 && 
b[54432] == 54432 && 
b[54433] == 54433 && 
b[54434] == 54434 && 
b[54435] == 54435 && 
b[54436] == 54436 && 
b[54437] == 54437 && 
b[54438] == 54438 && 
b[54439] == 54439 && 
b[54440] == 54440 && 
b[54441] == 54441 && 
b[54442] == 54442 && 
b[54443] == 54443 && 
b[54444] == 54444 && 
b[54445] == 54445 && 
b[54446] == 54446 && 
b[54447] == 54447 && 
b[54448] == 54448 && 
b[54449] == 54449 && 
b[54450] == 54450 && 
b[54451] == 54451 && 
b[54452] == 54452 && 
b[54453] == 54453 && 
b[54454] == 54454 && 
b[54455] == 54455 && 
b[54456] == 54456 && 
b[54457] == 54457 && 
b[54458] == 54458 && 
b[54459] == 54459 && 
b[54460] == 54460 && 
b[54461] == 54461 && 
b[54462] == 54462 && 
b[54463] == 54463 && 
b[54464] == 54464 && 
b[54465] == 54465 && 
b[54466] == 54466 && 
b[54467] == 54467 && 
b[54468] == 54468 && 
b[54469] == 54469 && 
b[54470] == 54470 && 
b[54471] == 54471 && 
b[54472] == 54472 && 
b[54473] == 54473 && 
b[54474] == 54474 && 
b[54475] == 54475 && 
b[54476] == 54476 && 
b[54477] == 54477 && 
b[54478] == 54478 && 
b[54479] == 54479 && 
b[54480] == 54480 && 
b[54481] == 54481 && 
b[54482] == 54482 && 
b[54483] == 54483 && 
b[54484] == 54484 && 
b[54485] == 54485 && 
b[54486] == 54486 && 
b[54487] == 54487 && 
b[54488] == 54488 && 
b[54489] == 54489 && 
b[54490] == 54490 && 
b[54491] == 54491 && 
b[54492] == 54492 && 
b[54493] == 54493 && 
b[54494] == 54494 && 
b[54495] == 54495 && 
b[54496] == 54496 && 
b[54497] == 54497 && 
b[54498] == 54498 && 
b[54499] == 54499 && 
b[54500] == 54500 && 
b[54501] == 54501 && 
b[54502] == 54502 && 
b[54503] == 54503 && 
b[54504] == 54504 && 
b[54505] == 54505 && 
b[54506] == 54506 && 
b[54507] == 54507 && 
b[54508] == 54508 && 
b[54509] == 54509 && 
b[54510] == 54510 && 
b[54511] == 54511 && 
b[54512] == 54512 && 
b[54513] == 54513 && 
b[54514] == 54514 && 
b[54515] == 54515 && 
b[54516] == 54516 && 
b[54517] == 54517 && 
b[54518] == 54518 && 
b[54519] == 54519 && 
b[54520] == 54520 && 
b[54521] == 54521 && 
b[54522] == 54522 && 
b[54523] == 54523 && 
b[54524] == 54524 && 
b[54525] == 54525 && 
b[54526] == 54526 && 
b[54527] == 54527 && 
b[54528] == 54528 && 
b[54529] == 54529 && 
b[54530] == 54530 && 
b[54531] == 54531 && 
b[54532] == 54532 && 
b[54533] == 54533 && 
b[54534] == 54534 && 
b[54535] == 54535 && 
b[54536] == 54536 && 
b[54537] == 54537 && 
b[54538] == 54538 && 
b[54539] == 54539 && 
b[54540] == 54540 && 
b[54541] == 54541 && 
b[54542] == 54542 && 
b[54543] == 54543 && 
b[54544] == 54544 && 
b[54545] == 54545 && 
b[54546] == 54546 && 
b[54547] == 54547 && 
b[54548] == 54548 && 
b[54549] == 54549 && 
b[54550] == 54550 && 
b[54551] == 54551 && 
b[54552] == 54552 && 
b[54553] == 54553 && 
b[54554] == 54554 && 
b[54555] == 54555 && 
b[54556] == 54556 && 
b[54557] == 54557 && 
b[54558] == 54558 && 
b[54559] == 54559 && 
b[54560] == 54560 && 
b[54561] == 54561 && 
b[54562] == 54562 && 
b[54563] == 54563 && 
b[54564] == 54564 && 
b[54565] == 54565 && 
b[54566] == 54566 && 
b[54567] == 54567 && 
b[54568] == 54568 && 
b[54569] == 54569 && 
b[54570] == 54570 && 
b[54571] == 54571 && 
b[54572] == 54572 && 
b[54573] == 54573 && 
b[54574] == 54574 && 
b[54575] == 54575 && 
b[54576] == 54576 && 
b[54577] == 54577 && 
b[54578] == 54578 && 
b[54579] == 54579 && 
b[54580] == 54580 && 
b[54581] == 54581 && 
b[54582] == 54582 && 
b[54583] == 54583 && 
b[54584] == 54584 && 
b[54585] == 54585 && 
b[54586] == 54586 && 
b[54587] == 54587 && 
b[54588] == 54588 && 
b[54589] == 54589 && 
b[54590] == 54590 && 
b[54591] == 54591 && 
b[54592] == 54592 && 
b[54593] == 54593 && 
b[54594] == 54594 && 
b[54595] == 54595 && 
b[54596] == 54596 && 
b[54597] == 54597 && 
b[54598] == 54598 && 
b[54599] == 54599 && 
b[54600] == 54600 && 
b[54601] == 54601 && 
b[54602] == 54602 && 
b[54603] == 54603 && 
b[54604] == 54604 && 
b[54605] == 54605 && 
b[54606] == 54606 && 
b[54607] == 54607 && 
b[54608] == 54608 && 
b[54609] == 54609 && 
b[54610] == 54610 && 
b[54611] == 54611 && 
b[54612] == 54612 && 
b[54613] == 54613 && 
b[54614] == 54614 && 
b[54615] == 54615 && 
b[54616] == 54616 && 
b[54617] == 54617 && 
b[54618] == 54618 && 
b[54619] == 54619 && 
b[54620] == 54620 && 
b[54621] == 54621 && 
b[54622] == 54622 && 
b[54623] == 54623 && 
b[54624] == 54624 && 
b[54625] == 54625 && 
b[54626] == 54626 && 
b[54627] == 54627 && 
b[54628] == 54628 && 
b[54629] == 54629 && 
b[54630] == 54630 && 
b[54631] == 54631 && 
b[54632] == 54632 && 
b[54633] == 54633 && 
b[54634] == 54634 && 
b[54635] == 54635 && 
b[54636] == 54636 && 
b[54637] == 54637 && 
b[54638] == 54638 && 
b[54639] == 54639 && 
b[54640] == 54640 && 
b[54641] == 54641 && 
b[54642] == 54642 && 
b[54643] == 54643 && 
b[54644] == 54644 && 
b[54645] == 54645 && 
b[54646] == 54646 && 
b[54647] == 54647 && 
b[54648] == 54648 && 
b[54649] == 54649 && 
b[54650] == 54650 && 
b[54651] == 54651 && 
b[54652] == 54652 && 
b[54653] == 54653 && 
b[54654] == 54654 && 
b[54655] == 54655 && 
b[54656] == 54656 && 
b[54657] == 54657 && 
b[54658] == 54658 && 
b[54659] == 54659 && 
b[54660] == 54660 && 
b[54661] == 54661 && 
b[54662] == 54662 && 
b[54663] == 54663 && 
b[54664] == 54664 && 
b[54665] == 54665 && 
b[54666] == 54666 && 
b[54667] == 54667 && 
b[54668] == 54668 && 
b[54669] == 54669 && 
b[54670] == 54670 && 
b[54671] == 54671 && 
b[54672] == 54672 && 
b[54673] == 54673 && 
b[54674] == 54674 && 
b[54675] == 54675 && 
b[54676] == 54676 && 
b[54677] == 54677 && 
b[54678] == 54678 && 
b[54679] == 54679 && 
b[54680] == 54680 && 
b[54681] == 54681 && 
b[54682] == 54682 && 
b[54683] == 54683 && 
b[54684] == 54684 && 
b[54685] == 54685 && 
b[54686] == 54686 && 
b[54687] == 54687 && 
b[54688] == 54688 && 
b[54689] == 54689 && 
b[54690] == 54690 && 
b[54691] == 54691 && 
b[54692] == 54692 && 
b[54693] == 54693 && 
b[54694] == 54694 && 
b[54695] == 54695 && 
b[54696] == 54696 && 
b[54697] == 54697 && 
b[54698] == 54698 && 
b[54699] == 54699 && 
b[54700] == 54700 && 
b[54701] == 54701 && 
b[54702] == 54702 && 
b[54703] == 54703 && 
b[54704] == 54704 && 
b[54705] == 54705 && 
b[54706] == 54706 && 
b[54707] == 54707 && 
b[54708] == 54708 && 
b[54709] == 54709 && 
b[54710] == 54710 && 
b[54711] == 54711 && 
b[54712] == 54712 && 
b[54713] == 54713 && 
b[54714] == 54714 && 
b[54715] == 54715 && 
b[54716] == 54716 && 
b[54717] == 54717 && 
b[54718] == 54718 && 
b[54719] == 54719 && 
b[54720] == 54720 && 
b[54721] == 54721 && 
b[54722] == 54722 && 
b[54723] == 54723 && 
b[54724] == 54724 && 
b[54725] == 54725 && 
b[54726] == 54726 && 
b[54727] == 54727 && 
b[54728] == 54728 && 
b[54729] == 54729 && 
b[54730] == 54730 && 
b[54731] == 54731 && 
b[54732] == 54732 && 
b[54733] == 54733 && 
b[54734] == 54734 && 
b[54735] == 54735 && 
b[54736] == 54736 && 
b[54737] == 54737 && 
b[54738] == 54738 && 
b[54739] == 54739 && 
b[54740] == 54740 && 
b[54741] == 54741 && 
b[54742] == 54742 && 
b[54743] == 54743 && 
b[54744] == 54744 && 
b[54745] == 54745 && 
b[54746] == 54746 && 
b[54747] == 54747 && 
b[54748] == 54748 && 
b[54749] == 54749 && 
b[54750] == 54750 && 
b[54751] == 54751 && 
b[54752] == 54752 && 
b[54753] == 54753 && 
b[54754] == 54754 && 
b[54755] == 54755 && 
b[54756] == 54756 && 
b[54757] == 54757 && 
b[54758] == 54758 && 
b[54759] == 54759 && 
b[54760] == 54760 && 
b[54761] == 54761 && 
b[54762] == 54762 && 
b[54763] == 54763 && 
b[54764] == 54764 && 
b[54765] == 54765 && 
b[54766] == 54766 && 
b[54767] == 54767 && 
b[54768] == 54768 && 
b[54769] == 54769 && 
b[54770] == 54770 && 
b[54771] == 54771 && 
b[54772] == 54772 && 
b[54773] == 54773 && 
b[54774] == 54774 && 
b[54775] == 54775 && 
b[54776] == 54776 && 
b[54777] == 54777 && 
b[54778] == 54778 && 
b[54779] == 54779 && 
b[54780] == 54780 && 
b[54781] == 54781 && 
b[54782] == 54782 && 
b[54783] == 54783 && 
b[54784] == 54784 && 
b[54785] == 54785 && 
b[54786] == 54786 && 
b[54787] == 54787 && 
b[54788] == 54788 && 
b[54789] == 54789 && 
b[54790] == 54790 && 
b[54791] == 54791 && 
b[54792] == 54792 && 
b[54793] == 54793 && 
b[54794] == 54794 && 
b[54795] == 54795 && 
b[54796] == 54796 && 
b[54797] == 54797 && 
b[54798] == 54798 && 
b[54799] == 54799 && 
b[54800] == 54800 && 
b[54801] == 54801 && 
b[54802] == 54802 && 
b[54803] == 54803 && 
b[54804] == 54804 && 
b[54805] == 54805 && 
b[54806] == 54806 && 
b[54807] == 54807 && 
b[54808] == 54808 && 
b[54809] == 54809 && 
b[54810] == 54810 && 
b[54811] == 54811 && 
b[54812] == 54812 && 
b[54813] == 54813 && 
b[54814] == 54814 && 
b[54815] == 54815 && 
b[54816] == 54816 && 
b[54817] == 54817 && 
b[54818] == 54818 && 
b[54819] == 54819 && 
b[54820] == 54820 && 
b[54821] == 54821 && 
b[54822] == 54822 && 
b[54823] == 54823 && 
b[54824] == 54824 && 
b[54825] == 54825 && 
b[54826] == 54826 && 
b[54827] == 54827 && 
b[54828] == 54828 && 
b[54829] == 54829 && 
b[54830] == 54830 && 
b[54831] == 54831 && 
b[54832] == 54832 && 
b[54833] == 54833 && 
b[54834] == 54834 && 
b[54835] == 54835 && 
b[54836] == 54836 && 
b[54837] == 54837 && 
b[54838] == 54838 && 
b[54839] == 54839 && 
b[54840] == 54840 && 
b[54841] == 54841 && 
b[54842] == 54842 && 
b[54843] == 54843 && 
b[54844] == 54844 && 
b[54845] == 54845 && 
b[54846] == 54846 && 
b[54847] == 54847 && 
b[54848] == 54848 && 
b[54849] == 54849 && 
b[54850] == 54850 && 
b[54851] == 54851 && 
b[54852] == 54852 && 
b[54853] == 54853 && 
b[54854] == 54854 && 
b[54855] == 54855 && 
b[54856] == 54856 && 
b[54857] == 54857 && 
b[54858] == 54858 && 
b[54859] == 54859 && 
b[54860] == 54860 && 
b[54861] == 54861 && 
b[54862] == 54862 && 
b[54863] == 54863 && 
b[54864] == 54864 && 
b[54865] == 54865 && 
b[54866] == 54866 && 
b[54867] == 54867 && 
b[54868] == 54868 && 
b[54869] == 54869 && 
b[54870] == 54870 && 
b[54871] == 54871 && 
b[54872] == 54872 && 
b[54873] == 54873 && 
b[54874] == 54874 && 
b[54875] == 54875 && 
b[54876] == 54876 && 
b[54877] == 54877 && 
b[54878] == 54878 && 
b[54879] == 54879 && 
b[54880] == 54880 && 
b[54881] == 54881 && 
b[54882] == 54882 && 
b[54883] == 54883 && 
b[54884] == 54884 && 
b[54885] == 54885 && 
b[54886] == 54886 && 
b[54887] == 54887 && 
b[54888] == 54888 && 
b[54889] == 54889 && 
b[54890] == 54890 && 
b[54891] == 54891 && 
b[54892] == 54892 && 
b[54893] == 54893 && 
b[54894] == 54894 && 
b[54895] == 54895 && 
b[54896] == 54896 && 
b[54897] == 54897 && 
b[54898] == 54898 && 
b[54899] == 54899 && 
b[54900] == 54900 && 
b[54901] == 54901 && 
b[54902] == 54902 && 
b[54903] == 54903 && 
b[54904] == 54904 && 
b[54905] == 54905 && 
b[54906] == 54906 && 
b[54907] == 54907 && 
b[54908] == 54908 && 
b[54909] == 54909 && 
b[54910] == 54910 && 
b[54911] == 54911 && 
b[54912] == 54912 && 
b[54913] == 54913 && 
b[54914] == 54914 && 
b[54915] == 54915 && 
b[54916] == 54916 && 
b[54917] == 54917 && 
b[54918] == 54918 && 
b[54919] == 54919 && 
b[54920] == 54920 && 
b[54921] == 54921 && 
b[54922] == 54922 && 
b[54923] == 54923 && 
b[54924] == 54924 && 
b[54925] == 54925 && 
b[54926] == 54926 && 
b[54927] == 54927 && 
b[54928] == 54928 && 
b[54929] == 54929 && 
b[54930] == 54930 && 
b[54931] == 54931 && 
b[54932] == 54932 && 
b[54933] == 54933 && 
b[54934] == 54934 && 
b[54935] == 54935 && 
b[54936] == 54936 && 
b[54937] == 54937 && 
b[54938] == 54938 && 
b[54939] == 54939 && 
b[54940] == 54940 && 
b[54941] == 54941 && 
b[54942] == 54942 && 
b[54943] == 54943 && 
b[54944] == 54944 && 
b[54945] == 54945 && 
b[54946] == 54946 && 
b[54947] == 54947 && 
b[54948] == 54948 && 
b[54949] == 54949 && 
b[54950] == 54950 && 
b[54951] == 54951 && 
b[54952] == 54952 && 
b[54953] == 54953 && 
b[54954] == 54954 && 
b[54955] == 54955 && 
b[54956] == 54956 && 
b[54957] == 54957 && 
b[54958] == 54958 && 
b[54959] == 54959 && 
b[54960] == 54960 && 
b[54961] == 54961 && 
b[54962] == 54962 && 
b[54963] == 54963 && 
b[54964] == 54964 && 
b[54965] == 54965 && 
b[54966] == 54966 && 
b[54967] == 54967 && 
b[54968] == 54968 && 
b[54969] == 54969 && 
b[54970] == 54970 && 
b[54971] == 54971 && 
b[54972] == 54972 && 
b[54973] == 54973 && 
b[54974] == 54974 && 
b[54975] == 54975 && 
b[54976] == 54976 && 
b[54977] == 54977 && 
b[54978] == 54978 && 
b[54979] == 54979 && 
b[54980] == 54980 && 
b[54981] == 54981 && 
b[54982] == 54982 && 
b[54983] == 54983 && 
b[54984] == 54984 && 
b[54985] == 54985 && 
b[54986] == 54986 && 
b[54987] == 54987 && 
b[54988] == 54988 && 
b[54989] == 54989 && 
b[54990] == 54990 && 
b[54991] == 54991 && 
b[54992] == 54992 && 
b[54993] == 54993 && 
b[54994] == 54994 && 
b[54995] == 54995 && 
b[54996] == 54996 && 
b[54997] == 54997 && 
b[54998] == 54998 && 
b[54999] == 54999 && 
b[55000] == 55000 && 
b[55001] == 55001 && 
b[55002] == 55002 && 
b[55003] == 55003 && 
b[55004] == 55004 && 
b[55005] == 55005 && 
b[55006] == 55006 && 
b[55007] == 55007 && 
b[55008] == 55008 && 
b[55009] == 55009 && 
b[55010] == 55010 && 
b[55011] == 55011 && 
b[55012] == 55012 && 
b[55013] == 55013 && 
b[55014] == 55014 && 
b[55015] == 55015 && 
b[55016] == 55016 && 
b[55017] == 55017 && 
b[55018] == 55018 && 
b[55019] == 55019 && 
b[55020] == 55020 && 
b[55021] == 55021 && 
b[55022] == 55022 && 
b[55023] == 55023 && 
b[55024] == 55024 && 
b[55025] == 55025 && 
b[55026] == 55026 && 
b[55027] == 55027 && 
b[55028] == 55028 && 
b[55029] == 55029 && 
b[55030] == 55030 && 
b[55031] == 55031 && 
b[55032] == 55032 && 
b[55033] == 55033 && 
b[55034] == 55034 && 
b[55035] == 55035 && 
b[55036] == 55036 && 
b[55037] == 55037 && 
b[55038] == 55038 && 
b[55039] == 55039 && 
b[55040] == 55040 && 
b[55041] == 55041 && 
b[55042] == 55042 && 
b[55043] == 55043 && 
b[55044] == 55044 && 
b[55045] == 55045 && 
b[55046] == 55046 && 
b[55047] == 55047 && 
b[55048] == 55048 && 
b[55049] == 55049 && 
b[55050] == 55050 && 
b[55051] == 55051 && 
b[55052] == 55052 && 
b[55053] == 55053 && 
b[55054] == 55054 && 
b[55055] == 55055 && 
b[55056] == 55056 && 
b[55057] == 55057 && 
b[55058] == 55058 && 
b[55059] == 55059 && 
b[55060] == 55060 && 
b[55061] == 55061 && 
b[55062] == 55062 && 
b[55063] == 55063 && 
b[55064] == 55064 && 
b[55065] == 55065 && 
b[55066] == 55066 && 
b[55067] == 55067 && 
b[55068] == 55068 && 
b[55069] == 55069 && 
b[55070] == 55070 && 
b[55071] == 55071 && 
b[55072] == 55072 && 
b[55073] == 55073 && 
b[55074] == 55074 && 
b[55075] == 55075 && 
b[55076] == 55076 && 
b[55077] == 55077 && 
b[55078] == 55078 && 
b[55079] == 55079 && 
b[55080] == 55080 && 
b[55081] == 55081 && 
b[55082] == 55082 && 
b[55083] == 55083 && 
b[55084] == 55084 && 
b[55085] == 55085 && 
b[55086] == 55086 && 
b[55087] == 55087 && 
b[55088] == 55088 && 
b[55089] == 55089 && 
b[55090] == 55090 && 
b[55091] == 55091 && 
b[55092] == 55092 && 
b[55093] == 55093 && 
b[55094] == 55094 && 
b[55095] == 55095 && 
b[55096] == 55096 && 
b[55097] == 55097 && 
b[55098] == 55098 && 
b[55099] == 55099 && 
b[55100] == 55100 && 
b[55101] == 55101 && 
b[55102] == 55102 && 
b[55103] == 55103 && 
b[55104] == 55104 && 
b[55105] == 55105 && 
b[55106] == 55106 && 
b[55107] == 55107 && 
b[55108] == 55108 && 
b[55109] == 55109 && 
b[55110] == 55110 && 
b[55111] == 55111 && 
b[55112] == 55112 && 
b[55113] == 55113 && 
b[55114] == 55114 && 
b[55115] == 55115 && 
b[55116] == 55116 && 
b[55117] == 55117 && 
b[55118] == 55118 && 
b[55119] == 55119 && 
b[55120] == 55120 && 
b[55121] == 55121 && 
b[55122] == 55122 && 
b[55123] == 55123 && 
b[55124] == 55124 && 
b[55125] == 55125 && 
b[55126] == 55126 && 
b[55127] == 55127 && 
b[55128] == 55128 && 
b[55129] == 55129 && 
b[55130] == 55130 && 
b[55131] == 55131 && 
b[55132] == 55132 && 
b[55133] == 55133 && 
b[55134] == 55134 && 
b[55135] == 55135 && 
b[55136] == 55136 && 
b[55137] == 55137 && 
b[55138] == 55138 && 
b[55139] == 55139 && 
b[55140] == 55140 && 
b[55141] == 55141 && 
b[55142] == 55142 && 
b[55143] == 55143 && 
b[55144] == 55144 && 
b[55145] == 55145 && 
b[55146] == 55146 && 
b[55147] == 55147 && 
b[55148] == 55148 && 
b[55149] == 55149 && 
b[55150] == 55150 && 
b[55151] == 55151 && 
b[55152] == 55152 && 
b[55153] == 55153 && 
b[55154] == 55154 && 
b[55155] == 55155 && 
b[55156] == 55156 && 
b[55157] == 55157 && 
b[55158] == 55158 && 
b[55159] == 55159 && 
b[55160] == 55160 && 
b[55161] == 55161 && 
b[55162] == 55162 && 
b[55163] == 55163 && 
b[55164] == 55164 && 
b[55165] == 55165 && 
b[55166] == 55166 && 
b[55167] == 55167 && 
b[55168] == 55168 && 
b[55169] == 55169 && 
b[55170] == 55170 && 
b[55171] == 55171 && 
b[55172] == 55172 && 
b[55173] == 55173 && 
b[55174] == 55174 && 
b[55175] == 55175 && 
b[55176] == 55176 && 
b[55177] == 55177 && 
b[55178] == 55178 && 
b[55179] == 55179 && 
b[55180] == 55180 && 
b[55181] == 55181 && 
b[55182] == 55182 && 
b[55183] == 55183 && 
b[55184] == 55184 && 
b[55185] == 55185 && 
b[55186] == 55186 && 
b[55187] == 55187 && 
b[55188] == 55188 && 
b[55189] == 55189 && 
b[55190] == 55190 && 
b[55191] == 55191 && 
b[55192] == 55192 && 
b[55193] == 55193 && 
b[55194] == 55194 && 
b[55195] == 55195 && 
b[55196] == 55196 && 
b[55197] == 55197 && 
b[55198] == 55198 && 
b[55199] == 55199 && 
b[55200] == 55200 && 
b[55201] == 55201 && 
b[55202] == 55202 && 
b[55203] == 55203 && 
b[55204] == 55204 && 
b[55205] == 55205 && 
b[55206] == 55206 && 
b[55207] == 55207 && 
b[55208] == 55208 && 
b[55209] == 55209 && 
b[55210] == 55210 && 
b[55211] == 55211 && 
b[55212] == 55212 && 
b[55213] == 55213 && 
b[55214] == 55214 && 
b[55215] == 55215 && 
b[55216] == 55216 && 
b[55217] == 55217 && 
b[55218] == 55218 && 
b[55219] == 55219 && 
b[55220] == 55220 && 
b[55221] == 55221 && 
b[55222] == 55222 && 
b[55223] == 55223 && 
b[55224] == 55224 && 
b[55225] == 55225 && 
b[55226] == 55226 && 
b[55227] == 55227 && 
b[55228] == 55228 && 
b[55229] == 55229 && 
b[55230] == 55230 && 
b[55231] == 55231 && 
b[55232] == 55232 && 
b[55233] == 55233 && 
b[55234] == 55234 && 
b[55235] == 55235 && 
b[55236] == 55236 && 
b[55237] == 55237 && 
b[55238] == 55238 && 
b[55239] == 55239 && 
b[55240] == 55240 && 
b[55241] == 55241 && 
b[55242] == 55242 && 
b[55243] == 55243 && 
b[55244] == 55244 && 
b[55245] == 55245 && 
b[55246] == 55246 && 
b[55247] == 55247 && 
b[55248] == 55248 && 
b[55249] == 55249 && 
b[55250] == 55250 && 
b[55251] == 55251 && 
b[55252] == 55252 && 
b[55253] == 55253 && 
b[55254] == 55254 && 
b[55255] == 55255 && 
b[55256] == 55256 && 
b[55257] == 55257 && 
b[55258] == 55258 && 
b[55259] == 55259 && 
b[55260] == 55260 && 
b[55261] == 55261 && 
b[55262] == 55262 && 
b[55263] == 55263 && 
b[55264] == 55264 && 
b[55265] == 55265 && 
b[55266] == 55266 && 
b[55267] == 55267 && 
b[55268] == 55268 && 
b[55269] == 55269 && 
b[55270] == 55270 && 
b[55271] == 55271 && 
b[55272] == 55272 && 
b[55273] == 55273 && 
b[55274] == 55274 && 
b[55275] == 55275 && 
b[55276] == 55276 && 
b[55277] == 55277 && 
b[55278] == 55278 && 
b[55279] == 55279 && 
b[55280] == 55280 && 
b[55281] == 55281 && 
b[55282] == 55282 && 
b[55283] == 55283 && 
b[55284] == 55284 && 
b[55285] == 55285 && 
b[55286] == 55286 && 
b[55287] == 55287 && 
b[55288] == 55288 && 
b[55289] == 55289 && 
b[55290] == 55290 && 
b[55291] == 55291 && 
b[55292] == 55292 && 
b[55293] == 55293 && 
b[55294] == 55294 && 
b[55295] == 55295 && 
b[55296] == 55296 && 
b[55297] == 55297 && 
b[55298] == 55298 && 
b[55299] == 55299 && 
b[55300] == 55300 && 
b[55301] == 55301 && 
b[55302] == 55302 && 
b[55303] == 55303 && 
b[55304] == 55304 && 
b[55305] == 55305 && 
b[55306] == 55306 && 
b[55307] == 55307 && 
b[55308] == 55308 && 
b[55309] == 55309 && 
b[55310] == 55310 && 
b[55311] == 55311 && 
b[55312] == 55312 && 
b[55313] == 55313 && 
b[55314] == 55314 && 
b[55315] == 55315 && 
b[55316] == 55316 && 
b[55317] == 55317 && 
b[55318] == 55318 && 
b[55319] == 55319 && 
b[55320] == 55320 && 
b[55321] == 55321 && 
b[55322] == 55322 && 
b[55323] == 55323 && 
b[55324] == 55324 && 
b[55325] == 55325 && 
b[55326] == 55326 && 
b[55327] == 55327 && 
b[55328] == 55328 && 
b[55329] == 55329 && 
b[55330] == 55330 && 
b[55331] == 55331 && 
b[55332] == 55332 && 
b[55333] == 55333 && 
b[55334] == 55334 && 
b[55335] == 55335 && 
b[55336] == 55336 && 
b[55337] == 55337 && 
b[55338] == 55338 && 
b[55339] == 55339 && 
b[55340] == 55340 && 
b[55341] == 55341 && 
b[55342] == 55342 && 
b[55343] == 55343 && 
b[55344] == 55344 && 
b[55345] == 55345 && 
b[55346] == 55346 && 
b[55347] == 55347 && 
b[55348] == 55348 && 
b[55349] == 55349 && 
b[55350] == 55350 && 
b[55351] == 55351 && 
b[55352] == 55352 && 
b[55353] == 55353 && 
b[55354] == 55354 && 
b[55355] == 55355 && 
b[55356] == 55356 && 
b[55357] == 55357 && 
b[55358] == 55358 && 
b[55359] == 55359 && 
b[55360] == 55360 && 
b[55361] == 55361 && 
b[55362] == 55362 && 
b[55363] == 55363 && 
b[55364] == 55364 && 
b[55365] == 55365 && 
b[55366] == 55366 && 
b[55367] == 55367 && 
b[55368] == 55368 && 
b[55369] == 55369 && 
b[55370] == 55370 && 
b[55371] == 55371 && 
b[55372] == 55372 && 
b[55373] == 55373 && 
b[55374] == 55374 && 
b[55375] == 55375 && 
b[55376] == 55376 && 
b[55377] == 55377 && 
b[55378] == 55378 && 
b[55379] == 55379 && 
b[55380] == 55380 && 
b[55381] == 55381 && 
b[55382] == 55382 && 
b[55383] == 55383 && 
b[55384] == 55384 && 
b[55385] == 55385 && 
b[55386] == 55386 && 
b[55387] == 55387 && 
b[55388] == 55388 && 
b[55389] == 55389 && 
b[55390] == 55390 && 
b[55391] == 55391 && 
b[55392] == 55392 && 
b[55393] == 55393 && 
b[55394] == 55394 && 
b[55395] == 55395 && 
b[55396] == 55396 && 
b[55397] == 55397 && 
b[55398] == 55398 && 
b[55399] == 55399 && 
b[55400] == 55400 && 
b[55401] == 55401 && 
b[55402] == 55402 && 
b[55403] == 55403 && 
b[55404] == 55404 && 
b[55405] == 55405 && 
b[55406] == 55406 && 
b[55407] == 55407 && 
b[55408] == 55408 && 
b[55409] == 55409 && 
b[55410] == 55410 && 
b[55411] == 55411 && 
b[55412] == 55412 && 
b[55413] == 55413 && 
b[55414] == 55414 && 
b[55415] == 55415 && 
b[55416] == 55416 && 
b[55417] == 55417 && 
b[55418] == 55418 && 
b[55419] == 55419 && 
b[55420] == 55420 && 
b[55421] == 55421 && 
b[55422] == 55422 && 
b[55423] == 55423 && 
b[55424] == 55424 && 
b[55425] == 55425 && 
b[55426] == 55426 && 
b[55427] == 55427 && 
b[55428] == 55428 && 
b[55429] == 55429 && 
b[55430] == 55430 && 
b[55431] == 55431 && 
b[55432] == 55432 && 
b[55433] == 55433 && 
b[55434] == 55434 && 
b[55435] == 55435 && 
b[55436] == 55436 && 
b[55437] == 55437 && 
b[55438] == 55438 && 
b[55439] == 55439 && 
b[55440] == 55440 && 
b[55441] == 55441 && 
b[55442] == 55442 && 
b[55443] == 55443 && 
b[55444] == 55444 && 
b[55445] == 55445 && 
b[55446] == 55446 && 
b[55447] == 55447 && 
b[55448] == 55448 && 
b[55449] == 55449 && 
b[55450] == 55450 && 
b[55451] == 55451 && 
b[55452] == 55452 && 
b[55453] == 55453 && 
b[55454] == 55454 && 
b[55455] == 55455 && 
b[55456] == 55456 && 
b[55457] == 55457 && 
b[55458] == 55458 && 
b[55459] == 55459 && 
b[55460] == 55460 && 
b[55461] == 55461 && 
b[55462] == 55462 && 
b[55463] == 55463 && 
b[55464] == 55464 && 
b[55465] == 55465 && 
b[55466] == 55466 && 
b[55467] == 55467 && 
b[55468] == 55468 && 
b[55469] == 55469 && 
b[55470] == 55470 && 
b[55471] == 55471 && 
b[55472] == 55472 && 
b[55473] == 55473 && 
b[55474] == 55474 && 
b[55475] == 55475 && 
b[55476] == 55476 && 
b[55477] == 55477 && 
b[55478] == 55478 && 
b[55479] == 55479 && 
b[55480] == 55480 && 
b[55481] == 55481 && 
b[55482] == 55482 && 
b[55483] == 55483 && 
b[55484] == 55484 && 
b[55485] == 55485 && 
b[55486] == 55486 && 
b[55487] == 55487 && 
b[55488] == 55488 && 
b[55489] == 55489 && 
b[55490] == 55490 && 
b[55491] == 55491 && 
b[55492] == 55492 && 
b[55493] == 55493 && 
b[55494] == 55494 && 
b[55495] == 55495 && 
b[55496] == 55496 && 
b[55497] == 55497 && 
b[55498] == 55498 && 
b[55499] == 55499 && 
b[55500] == 55500 && 
b[55501] == 55501 && 
b[55502] == 55502 && 
b[55503] == 55503 && 
b[55504] == 55504 && 
b[55505] == 55505 && 
b[55506] == 55506 && 
b[55507] == 55507 && 
b[55508] == 55508 && 
b[55509] == 55509 && 
b[55510] == 55510 && 
b[55511] == 55511 && 
b[55512] == 55512 && 
b[55513] == 55513 && 
b[55514] == 55514 && 
b[55515] == 55515 && 
b[55516] == 55516 && 
b[55517] == 55517 && 
b[55518] == 55518 && 
b[55519] == 55519 && 
b[55520] == 55520 && 
b[55521] == 55521 && 
b[55522] == 55522 && 
b[55523] == 55523 && 
b[55524] == 55524 && 
b[55525] == 55525 && 
b[55526] == 55526 && 
b[55527] == 55527 && 
b[55528] == 55528 && 
b[55529] == 55529 && 
b[55530] == 55530 && 
b[55531] == 55531 && 
b[55532] == 55532 && 
b[55533] == 55533 && 
b[55534] == 55534 && 
b[55535] == 55535 && 
b[55536] == 55536 && 
b[55537] == 55537 && 
b[55538] == 55538 && 
b[55539] == 55539 && 
b[55540] == 55540 && 
b[55541] == 55541 && 
b[55542] == 55542 && 
b[55543] == 55543 && 
b[55544] == 55544 && 
b[55545] == 55545 && 
b[55546] == 55546 && 
b[55547] == 55547 && 
b[55548] == 55548 && 
b[55549] == 55549 && 
b[55550] == 55550 && 
b[55551] == 55551 && 
b[55552] == 55552 && 
b[55553] == 55553 && 
b[55554] == 55554 && 
b[55555] == 55555 && 
b[55556] == 55556 && 
b[55557] == 55557 && 
b[55558] == 55558 && 
b[55559] == 55559 && 
b[55560] == 55560 && 
b[55561] == 55561 && 
b[55562] == 55562 && 
b[55563] == 55563 && 
b[55564] == 55564 && 
b[55565] == 55565 && 
b[55566] == 55566 && 
b[55567] == 55567 && 
b[55568] == 55568 && 
b[55569] == 55569 && 
b[55570] == 55570 && 
b[55571] == 55571 && 
b[55572] == 55572 && 
b[55573] == 55573 && 
b[55574] == 55574 && 
b[55575] == 55575 && 
b[55576] == 55576 && 
b[55577] == 55577 && 
b[55578] == 55578 && 
b[55579] == 55579 && 
b[55580] == 55580 && 
b[55581] == 55581 && 
b[55582] == 55582 && 
b[55583] == 55583 && 
b[55584] == 55584 && 
b[55585] == 55585 && 
b[55586] == 55586 && 
b[55587] == 55587 && 
b[55588] == 55588 && 
b[55589] == 55589 && 
b[55590] == 55590 && 
b[55591] == 55591 && 
b[55592] == 55592 && 
b[55593] == 55593 && 
b[55594] == 55594 && 
b[55595] == 55595 && 
b[55596] == 55596 && 
b[55597] == 55597 && 
b[55598] == 55598 && 
b[55599] == 55599 && 
b[55600] == 55600 && 
b[55601] == 55601 && 
b[55602] == 55602 && 
b[55603] == 55603 && 
b[55604] == 55604 && 
b[55605] == 55605 && 
b[55606] == 55606 && 
b[55607] == 55607 && 
b[55608] == 55608 && 
b[55609] == 55609 && 
b[55610] == 55610 && 
b[55611] == 55611 && 
b[55612] == 55612 && 
b[55613] == 55613 && 
b[55614] == 55614 && 
b[55615] == 55615 && 
b[55616] == 55616 && 
b[55617] == 55617 && 
b[55618] == 55618 && 
b[55619] == 55619 && 
b[55620] == 55620 && 
b[55621] == 55621 && 
b[55622] == 55622 && 
b[55623] == 55623 && 
b[55624] == 55624 && 
b[55625] == 55625 && 
b[55626] == 55626 && 
b[55627] == 55627 && 
b[55628] == 55628 && 
b[55629] == 55629 && 
b[55630] == 55630 && 
b[55631] == 55631 && 
b[55632] == 55632 && 
b[55633] == 55633 && 
b[55634] == 55634 && 
b[55635] == 55635 && 
b[55636] == 55636 && 
b[55637] == 55637 && 
b[55638] == 55638 && 
b[55639] == 55639 && 
b[55640] == 55640 && 
b[55641] == 55641 && 
b[55642] == 55642 && 
b[55643] == 55643 && 
b[55644] == 55644 && 
b[55645] == 55645 && 
b[55646] == 55646 && 
b[55647] == 55647 && 
b[55648] == 55648 && 
b[55649] == 55649 && 
b[55650] == 55650 && 
b[55651] == 55651 && 
b[55652] == 55652 && 
b[55653] == 55653 && 
b[55654] == 55654 && 
b[55655] == 55655 && 
b[55656] == 55656 && 
b[55657] == 55657 && 
b[55658] == 55658 && 
b[55659] == 55659 && 
b[55660] == 55660 && 
b[55661] == 55661 && 
b[55662] == 55662 && 
b[55663] == 55663 && 
b[55664] == 55664 && 
b[55665] == 55665 && 
b[55666] == 55666 && 
b[55667] == 55667 && 
b[55668] == 55668 && 
b[55669] == 55669 && 
b[55670] == 55670 && 
b[55671] == 55671 && 
b[55672] == 55672 && 
b[55673] == 55673 && 
b[55674] == 55674 && 
b[55675] == 55675 && 
b[55676] == 55676 && 
b[55677] == 55677 && 
b[55678] == 55678 && 
b[55679] == 55679 && 
b[55680] == 55680 && 
b[55681] == 55681 && 
b[55682] == 55682 && 
b[55683] == 55683 && 
b[55684] == 55684 && 
b[55685] == 55685 && 
b[55686] == 55686 && 
b[55687] == 55687 && 
b[55688] == 55688 && 
b[55689] == 55689 && 
b[55690] == 55690 && 
b[55691] == 55691 && 
b[55692] == 55692 && 
b[55693] == 55693 && 
b[55694] == 55694 && 
b[55695] == 55695 && 
b[55696] == 55696 && 
b[55697] == 55697 && 
b[55698] == 55698 && 
b[55699] == 55699 && 
b[55700] == 55700 && 
b[55701] == 55701 && 
b[55702] == 55702 && 
b[55703] == 55703 && 
b[55704] == 55704 && 
b[55705] == 55705 && 
b[55706] == 55706 && 
b[55707] == 55707 && 
b[55708] == 55708 && 
b[55709] == 55709 && 
b[55710] == 55710 && 
b[55711] == 55711 && 
b[55712] == 55712 && 
b[55713] == 55713 && 
b[55714] == 55714 && 
b[55715] == 55715 && 
b[55716] == 55716 && 
b[55717] == 55717 && 
b[55718] == 55718 && 
b[55719] == 55719 && 
b[55720] == 55720 && 
b[55721] == 55721 && 
b[55722] == 55722 && 
b[55723] == 55723 && 
b[55724] == 55724 && 
b[55725] == 55725 && 
b[55726] == 55726 && 
b[55727] == 55727 && 
b[55728] == 55728 && 
b[55729] == 55729 && 
b[55730] == 55730 && 
b[55731] == 55731 && 
b[55732] == 55732 && 
b[55733] == 55733 && 
b[55734] == 55734 && 
b[55735] == 55735 && 
b[55736] == 55736 && 
b[55737] == 55737 && 
b[55738] == 55738 && 
b[55739] == 55739 && 
b[55740] == 55740 && 
b[55741] == 55741 && 
b[55742] == 55742 && 
b[55743] == 55743 && 
b[55744] == 55744 && 
b[55745] == 55745 && 
b[55746] == 55746 && 
b[55747] == 55747 && 
b[55748] == 55748 && 
b[55749] == 55749 && 
b[55750] == 55750 && 
b[55751] == 55751 && 
b[55752] == 55752 && 
b[55753] == 55753 && 
b[55754] == 55754 && 
b[55755] == 55755 && 
b[55756] == 55756 && 
b[55757] == 55757 && 
b[55758] == 55758 && 
b[55759] == 55759 && 
b[55760] == 55760 && 
b[55761] == 55761 && 
b[55762] == 55762 && 
b[55763] == 55763 && 
b[55764] == 55764 && 
b[55765] == 55765 && 
b[55766] == 55766 && 
b[55767] == 55767 && 
b[55768] == 55768 && 
b[55769] == 55769 && 
b[55770] == 55770 && 
b[55771] == 55771 && 
b[55772] == 55772 && 
b[55773] == 55773 && 
b[55774] == 55774 && 
b[55775] == 55775 && 
b[55776] == 55776 && 
b[55777] == 55777 && 
b[55778] == 55778 && 
b[55779] == 55779 && 
b[55780] == 55780 && 
b[55781] == 55781 && 
b[55782] == 55782 && 
b[55783] == 55783 && 
b[55784] == 55784 && 
b[55785] == 55785 && 
b[55786] == 55786 && 
b[55787] == 55787 && 
b[55788] == 55788 && 
b[55789] == 55789 && 
b[55790] == 55790 && 
b[55791] == 55791 && 
b[55792] == 55792 && 
b[55793] == 55793 && 
b[55794] == 55794 && 
b[55795] == 55795 && 
b[55796] == 55796 && 
b[55797] == 55797 && 
b[55798] == 55798 && 
b[55799] == 55799 && 
b[55800] == 55800 && 
b[55801] == 55801 && 
b[55802] == 55802 && 
b[55803] == 55803 && 
b[55804] == 55804 && 
b[55805] == 55805 && 
b[55806] == 55806 && 
b[55807] == 55807 && 
b[55808] == 55808 && 
b[55809] == 55809 && 
b[55810] == 55810 && 
b[55811] == 55811 && 
b[55812] == 55812 && 
b[55813] == 55813 && 
b[55814] == 55814 && 
b[55815] == 55815 && 
b[55816] == 55816 && 
b[55817] == 55817 && 
b[55818] == 55818 && 
b[55819] == 55819 && 
b[55820] == 55820 && 
b[55821] == 55821 && 
b[55822] == 55822 && 
b[55823] == 55823 && 
b[55824] == 55824 && 
b[55825] == 55825 && 
b[55826] == 55826 && 
b[55827] == 55827 && 
b[55828] == 55828 && 
b[55829] == 55829 && 
b[55830] == 55830 && 
b[55831] == 55831 && 
b[55832] == 55832 && 
b[55833] == 55833 && 
b[55834] == 55834 && 
b[55835] == 55835 && 
b[55836] == 55836 && 
b[55837] == 55837 && 
b[55838] == 55838 && 
b[55839] == 55839 && 
b[55840] == 55840 && 
b[55841] == 55841 && 
b[55842] == 55842 && 
b[55843] == 55843 && 
b[55844] == 55844 && 
b[55845] == 55845 && 
b[55846] == 55846 && 
b[55847] == 55847 && 
b[55848] == 55848 && 
b[55849] == 55849 && 
b[55850] == 55850 && 
b[55851] == 55851 && 
b[55852] == 55852 && 
b[55853] == 55853 && 
b[55854] == 55854 && 
b[55855] == 55855 && 
b[55856] == 55856 && 
b[55857] == 55857 && 
b[55858] == 55858 && 
b[55859] == 55859 && 
b[55860] == 55860 && 
b[55861] == 55861 && 
b[55862] == 55862 && 
b[55863] == 55863 && 
b[55864] == 55864 && 
b[55865] == 55865 && 
b[55866] == 55866 && 
b[55867] == 55867 && 
b[55868] == 55868 && 
b[55869] == 55869 && 
b[55870] == 55870 && 
b[55871] == 55871 && 
b[55872] == 55872 && 
b[55873] == 55873 && 
b[55874] == 55874 && 
b[55875] == 55875 && 
b[55876] == 55876 && 
b[55877] == 55877 && 
b[55878] == 55878 && 
b[55879] == 55879 && 
b[55880] == 55880 && 
b[55881] == 55881 && 
b[55882] == 55882 && 
b[55883] == 55883 && 
b[55884] == 55884 && 
b[55885] == 55885 && 
b[55886] == 55886 && 
b[55887] == 55887 && 
b[55888] == 55888 && 
b[55889] == 55889 && 
b[55890] == 55890 && 
b[55891] == 55891 && 
b[55892] == 55892 && 
b[55893] == 55893 && 
b[55894] == 55894 && 
b[55895] == 55895 && 
b[55896] == 55896 && 
b[55897] == 55897 && 
b[55898] == 55898 && 
b[55899] == 55899 && 
b[55900] == 55900 && 
b[55901] == 55901 && 
b[55902] == 55902 && 
b[55903] == 55903 && 
b[55904] == 55904 && 
b[55905] == 55905 && 
b[55906] == 55906 && 
b[55907] == 55907 && 
b[55908] == 55908 && 
b[55909] == 55909 && 
b[55910] == 55910 && 
b[55911] == 55911 && 
b[55912] == 55912 && 
b[55913] == 55913 && 
b[55914] == 55914 && 
b[55915] == 55915 && 
b[55916] == 55916 && 
b[55917] == 55917 && 
b[55918] == 55918 && 
b[55919] == 55919 && 
b[55920] == 55920 && 
b[55921] == 55921 && 
b[55922] == 55922 && 
b[55923] == 55923 && 
b[55924] == 55924 && 
b[55925] == 55925 && 
b[55926] == 55926 && 
b[55927] == 55927 && 
b[55928] == 55928 && 
b[55929] == 55929 && 
b[55930] == 55930 && 
b[55931] == 55931 && 
b[55932] == 55932 && 
b[55933] == 55933 && 
b[55934] == 55934 && 
b[55935] == 55935 && 
b[55936] == 55936 && 
b[55937] == 55937 && 
b[55938] == 55938 && 
b[55939] == 55939 && 
b[55940] == 55940 && 
b[55941] == 55941 && 
b[55942] == 55942 && 
b[55943] == 55943 && 
b[55944] == 55944 && 
b[55945] == 55945 && 
b[55946] == 55946 && 
b[55947] == 55947 && 
b[55948] == 55948 && 
b[55949] == 55949 && 
b[55950] == 55950 && 
b[55951] == 55951 && 
b[55952] == 55952 && 
b[55953] == 55953 && 
b[55954] == 55954 && 
b[55955] == 55955 && 
b[55956] == 55956 && 
b[55957] == 55957 && 
b[55958] == 55958 && 
b[55959] == 55959 && 
b[55960] == 55960 && 
b[55961] == 55961 && 
b[55962] == 55962 && 
b[55963] == 55963 && 
b[55964] == 55964 && 
b[55965] == 55965 && 
b[55966] == 55966 && 
b[55967] == 55967 && 
b[55968] == 55968 && 
b[55969] == 55969 && 
b[55970] == 55970 && 
b[55971] == 55971 && 
b[55972] == 55972 && 
b[55973] == 55973 && 
b[55974] == 55974 && 
b[55975] == 55975 && 
b[55976] == 55976 && 
b[55977] == 55977 && 
b[55978] == 55978 && 
b[55979] == 55979 && 
b[55980] == 55980 && 
b[55981] == 55981 && 
b[55982] == 55982 && 
b[55983] == 55983 && 
b[55984] == 55984 && 
b[55985] == 55985 && 
b[55986] == 55986 && 
b[55987] == 55987 && 
b[55988] == 55988 && 
b[55989] == 55989 && 
b[55990] == 55990 && 
b[55991] == 55991 && 
b[55992] == 55992 && 
b[55993] == 55993 && 
b[55994] == 55994 && 
b[55995] == 55995 && 
b[55996] == 55996 && 
b[55997] == 55997 && 
b[55998] == 55998 && 
b[55999] == 55999 && 
b[56000] == 56000 && 
b[56001] == 56001 && 
b[56002] == 56002 && 
b[56003] == 56003 && 
b[56004] == 56004 && 
b[56005] == 56005 && 
b[56006] == 56006 && 
b[56007] == 56007 && 
b[56008] == 56008 && 
b[56009] == 56009 && 
b[56010] == 56010 && 
b[56011] == 56011 && 
b[56012] == 56012 && 
b[56013] == 56013 && 
b[56014] == 56014 && 
b[56015] == 56015 && 
b[56016] == 56016 && 
b[56017] == 56017 && 
b[56018] == 56018 && 
b[56019] == 56019 && 
b[56020] == 56020 && 
b[56021] == 56021 && 
b[56022] == 56022 && 
b[56023] == 56023 && 
b[56024] == 56024 && 
b[56025] == 56025 && 
b[56026] == 56026 && 
b[56027] == 56027 && 
b[56028] == 56028 && 
b[56029] == 56029 && 
b[56030] == 56030 && 
b[56031] == 56031 && 
b[56032] == 56032 && 
b[56033] == 56033 && 
b[56034] == 56034 && 
b[56035] == 56035 && 
b[56036] == 56036 && 
b[56037] == 56037 && 
b[56038] == 56038 && 
b[56039] == 56039 && 
b[56040] == 56040 && 
b[56041] == 56041 && 
b[56042] == 56042 && 
b[56043] == 56043 && 
b[56044] == 56044 && 
b[56045] == 56045 && 
b[56046] == 56046 && 
b[56047] == 56047 && 
b[56048] == 56048 && 
b[56049] == 56049 && 
b[56050] == 56050 && 
b[56051] == 56051 && 
b[56052] == 56052 && 
b[56053] == 56053 && 
b[56054] == 56054 && 
b[56055] == 56055 && 
b[56056] == 56056 && 
b[56057] == 56057 && 
b[56058] == 56058 && 
b[56059] == 56059 && 
b[56060] == 56060 && 
b[56061] == 56061 && 
b[56062] == 56062 && 
b[56063] == 56063 && 
b[56064] == 56064 && 
b[56065] == 56065 && 
b[56066] == 56066 && 
b[56067] == 56067 && 
b[56068] == 56068 && 
b[56069] == 56069 && 
b[56070] == 56070 && 
b[56071] == 56071 && 
b[56072] == 56072 && 
b[56073] == 56073 && 
b[56074] == 56074 && 
b[56075] == 56075 && 
b[56076] == 56076 && 
b[56077] == 56077 && 
b[56078] == 56078 && 
b[56079] == 56079 && 
b[56080] == 56080 && 
b[56081] == 56081 && 
b[56082] == 56082 && 
b[56083] == 56083 && 
b[56084] == 56084 && 
b[56085] == 56085 && 
b[56086] == 56086 && 
b[56087] == 56087 && 
b[56088] == 56088 && 
b[56089] == 56089 && 
b[56090] == 56090 && 
b[56091] == 56091 && 
b[56092] == 56092 && 
b[56093] == 56093 && 
b[56094] == 56094 && 
b[56095] == 56095 && 
b[56096] == 56096 && 
b[56097] == 56097 && 
b[56098] == 56098 && 
b[56099] == 56099 && 
b[56100] == 56100 && 
b[56101] == 56101 && 
b[56102] == 56102 && 
b[56103] == 56103 && 
b[56104] == 56104 && 
b[56105] == 56105 && 
b[56106] == 56106 && 
b[56107] == 56107 && 
b[56108] == 56108 && 
b[56109] == 56109 && 
b[56110] == 56110 && 
b[56111] == 56111 && 
b[56112] == 56112 && 
b[56113] == 56113 && 
b[56114] == 56114 && 
b[56115] == 56115 && 
b[56116] == 56116 && 
b[56117] == 56117 && 
b[56118] == 56118 && 
b[56119] == 56119 && 
b[56120] == 56120 && 
b[56121] == 56121 && 
b[56122] == 56122 && 
b[56123] == 56123 && 
b[56124] == 56124 && 
b[56125] == 56125 && 
b[56126] == 56126 && 
b[56127] == 56127 && 
b[56128] == 56128 && 
b[56129] == 56129 && 
b[56130] == 56130 && 
b[56131] == 56131 && 
b[56132] == 56132 && 
b[56133] == 56133 && 
b[56134] == 56134 && 
b[56135] == 56135 && 
b[56136] == 56136 && 
b[56137] == 56137 && 
b[56138] == 56138 && 
b[56139] == 56139 && 
b[56140] == 56140 && 
b[56141] == 56141 && 
b[56142] == 56142 && 
b[56143] == 56143 && 
b[56144] == 56144 && 
b[56145] == 56145 && 
b[56146] == 56146 && 
b[56147] == 56147 && 
b[56148] == 56148 && 
b[56149] == 56149 && 
b[56150] == 56150 && 
b[56151] == 56151 && 
b[56152] == 56152 && 
b[56153] == 56153 && 
b[56154] == 56154 && 
b[56155] == 56155 && 
b[56156] == 56156 && 
b[56157] == 56157 && 
b[56158] == 56158 && 
b[56159] == 56159 && 
b[56160] == 56160 && 
b[56161] == 56161 && 
b[56162] == 56162 && 
b[56163] == 56163 && 
b[56164] == 56164 && 
b[56165] == 56165 && 
b[56166] == 56166 && 
b[56167] == 56167 && 
b[56168] == 56168 && 
b[56169] == 56169 && 
b[56170] == 56170 && 
b[56171] == 56171 && 
b[56172] == 56172 && 
b[56173] == 56173 && 
b[56174] == 56174 && 
b[56175] == 56175 && 
b[56176] == 56176 && 
b[56177] == 56177 && 
b[56178] == 56178 && 
b[56179] == 56179 && 
b[56180] == 56180 && 
b[56181] == 56181 && 
b[56182] == 56182 && 
b[56183] == 56183 && 
b[56184] == 56184 && 
b[56185] == 56185 && 
b[56186] == 56186 && 
b[56187] == 56187 && 
b[56188] == 56188 && 
b[56189] == 56189 && 
b[56190] == 56190 && 
b[56191] == 56191 && 
b[56192] == 56192 && 
b[56193] == 56193 && 
b[56194] == 56194 && 
b[56195] == 56195 && 
b[56196] == 56196 && 
b[56197] == 56197 && 
b[56198] == 56198 && 
b[56199] == 56199 && 
b[56200] == 56200 && 
b[56201] == 56201 && 
b[56202] == 56202 && 
b[56203] == 56203 && 
b[56204] == 56204 && 
b[56205] == 56205 && 
b[56206] == 56206 && 
b[56207] == 56207 && 
b[56208] == 56208 && 
b[56209] == 56209 && 
b[56210] == 56210 && 
b[56211] == 56211 && 
b[56212] == 56212 && 
b[56213] == 56213 && 
b[56214] == 56214 && 
b[56215] == 56215 && 
b[56216] == 56216 && 
b[56217] == 56217 && 
b[56218] == 56218 && 
b[56219] == 56219 && 
b[56220] == 56220 && 
b[56221] == 56221 && 
b[56222] == 56222 && 
b[56223] == 56223 && 
b[56224] == 56224 && 
b[56225] == 56225 && 
b[56226] == 56226 && 
b[56227] == 56227 && 
b[56228] == 56228 && 
b[56229] == 56229 && 
b[56230] == 56230 && 
b[56231] == 56231 && 
b[56232] == 56232 && 
b[56233] == 56233 && 
b[56234] == 56234 && 
b[56235] == 56235 && 
b[56236] == 56236 && 
b[56237] == 56237 && 
b[56238] == 56238 && 
b[56239] == 56239 && 
b[56240] == 56240 && 
b[56241] == 56241 && 
b[56242] == 56242 && 
b[56243] == 56243 && 
b[56244] == 56244 && 
b[56245] == 56245 && 
b[56246] == 56246 && 
b[56247] == 56247 && 
b[56248] == 56248 && 
b[56249] == 56249 && 
b[56250] == 56250 && 
b[56251] == 56251 && 
b[56252] == 56252 && 
b[56253] == 56253 && 
b[56254] == 56254 && 
b[56255] == 56255 && 
b[56256] == 56256 && 
b[56257] == 56257 && 
b[56258] == 56258 && 
b[56259] == 56259 && 
b[56260] == 56260 && 
b[56261] == 56261 && 
b[56262] == 56262 && 
b[56263] == 56263 && 
b[56264] == 56264 && 
b[56265] == 56265 && 
b[56266] == 56266 && 
b[56267] == 56267 && 
b[56268] == 56268 && 
b[56269] == 56269 && 
b[56270] == 56270 && 
b[56271] == 56271 && 
b[56272] == 56272 && 
b[56273] == 56273 && 
b[56274] == 56274 && 
b[56275] == 56275 && 
b[56276] == 56276 && 
b[56277] == 56277 && 
b[56278] == 56278 && 
b[56279] == 56279 && 
b[56280] == 56280 && 
b[56281] == 56281 && 
b[56282] == 56282 && 
b[56283] == 56283 && 
b[56284] == 56284 && 
b[56285] == 56285 && 
b[56286] == 56286 && 
b[56287] == 56287 && 
b[56288] == 56288 && 
b[56289] == 56289 && 
b[56290] == 56290 && 
b[56291] == 56291 && 
b[56292] == 56292 && 
b[56293] == 56293 && 
b[56294] == 56294 && 
b[56295] == 56295 && 
b[56296] == 56296 && 
b[56297] == 56297 && 
b[56298] == 56298 && 
b[56299] == 56299 && 
b[56300] == 56300 && 
b[56301] == 56301 && 
b[56302] == 56302 && 
b[56303] == 56303 && 
b[56304] == 56304 && 
b[56305] == 56305 && 
b[56306] == 56306 && 
b[56307] == 56307 && 
b[56308] == 56308 && 
b[56309] == 56309 && 
b[56310] == 56310 && 
b[56311] == 56311 && 
b[56312] == 56312 && 
b[56313] == 56313 && 
b[56314] == 56314 && 
b[56315] == 56315 && 
b[56316] == 56316 && 
b[56317] == 56317 && 
b[56318] == 56318 && 
b[56319] == 56319 && 
b[56320] == 56320 && 
b[56321] == 56321 && 
b[56322] == 56322 && 
b[56323] == 56323 && 
b[56324] == 56324 && 
b[56325] == 56325 && 
b[56326] == 56326 && 
b[56327] == 56327 && 
b[56328] == 56328 && 
b[56329] == 56329 && 
b[56330] == 56330 && 
b[56331] == 56331 && 
b[56332] == 56332 && 
b[56333] == 56333 && 
b[56334] == 56334 && 
b[56335] == 56335 && 
b[56336] == 56336 && 
b[56337] == 56337 && 
b[56338] == 56338 && 
b[56339] == 56339 && 
b[56340] == 56340 && 
b[56341] == 56341 && 
b[56342] == 56342 && 
b[56343] == 56343 && 
b[56344] == 56344 && 
b[56345] == 56345 && 
b[56346] == 56346 && 
b[56347] == 56347 && 
b[56348] == 56348 && 
b[56349] == 56349 && 
b[56350] == 56350 && 
b[56351] == 56351 && 
b[56352] == 56352 && 
b[56353] == 56353 && 
b[56354] == 56354 && 
b[56355] == 56355 && 
b[56356] == 56356 && 
b[56357] == 56357 && 
b[56358] == 56358 && 
b[56359] == 56359 && 
b[56360] == 56360 && 
b[56361] == 56361 && 
b[56362] == 56362 && 
b[56363] == 56363 && 
b[56364] == 56364 && 
b[56365] == 56365 && 
b[56366] == 56366 && 
b[56367] == 56367 && 
b[56368] == 56368 && 
b[56369] == 56369 && 
b[56370] == 56370 && 
b[56371] == 56371 && 
b[56372] == 56372 && 
b[56373] == 56373 && 
b[56374] == 56374 && 
b[56375] == 56375 && 
b[56376] == 56376 && 
b[56377] == 56377 && 
b[56378] == 56378 && 
b[56379] == 56379 && 
b[56380] == 56380 && 
b[56381] == 56381 && 
b[56382] == 56382 && 
b[56383] == 56383 && 
b[56384] == 56384 && 
b[56385] == 56385 && 
b[56386] == 56386 && 
b[56387] == 56387 && 
b[56388] == 56388 && 
b[56389] == 56389 && 
b[56390] == 56390 && 
b[56391] == 56391 && 
b[56392] == 56392 && 
b[56393] == 56393 && 
b[56394] == 56394 && 
b[56395] == 56395 && 
b[56396] == 56396 && 
b[56397] == 56397 && 
b[56398] == 56398 && 
b[56399] == 56399 && 
b[56400] == 56400 && 
b[56401] == 56401 && 
b[56402] == 56402 && 
b[56403] == 56403 && 
b[56404] == 56404 && 
b[56405] == 56405 && 
b[56406] == 56406 && 
b[56407] == 56407 && 
b[56408] == 56408 && 
b[56409] == 56409 && 
b[56410] == 56410 && 
b[56411] == 56411 && 
b[56412] == 56412 && 
b[56413] == 56413 && 
b[56414] == 56414 && 
b[56415] == 56415 && 
b[56416] == 56416 && 
b[56417] == 56417 && 
b[56418] == 56418 && 
b[56419] == 56419 && 
b[56420] == 56420 && 
b[56421] == 56421 && 
b[56422] == 56422 && 
b[56423] == 56423 && 
b[56424] == 56424 && 
b[56425] == 56425 && 
b[56426] == 56426 && 
b[56427] == 56427 && 
b[56428] == 56428 && 
b[56429] == 56429 && 
b[56430] == 56430 && 
b[56431] == 56431 && 
b[56432] == 56432 && 
b[56433] == 56433 && 
b[56434] == 56434 && 
b[56435] == 56435 && 
b[56436] == 56436 && 
b[56437] == 56437 && 
b[56438] == 56438 && 
b[56439] == 56439 && 
b[56440] == 56440 && 
b[56441] == 56441 && 
b[56442] == 56442 && 
b[56443] == 56443 && 
b[56444] == 56444 && 
b[56445] == 56445 && 
b[56446] == 56446 && 
b[56447] == 56447 && 
b[56448] == 56448 && 
b[56449] == 56449 && 
b[56450] == 56450 && 
b[56451] == 56451 && 
b[56452] == 56452 && 
b[56453] == 56453 && 
b[56454] == 56454 && 
b[56455] == 56455 && 
b[56456] == 56456 && 
b[56457] == 56457 && 
b[56458] == 56458 && 
b[56459] == 56459 && 
b[56460] == 56460 && 
b[56461] == 56461 && 
b[56462] == 56462 && 
b[56463] == 56463 && 
b[56464] == 56464 && 
b[56465] == 56465 && 
b[56466] == 56466 && 
b[56467] == 56467 && 
b[56468] == 56468 && 
b[56469] == 56469 && 
b[56470] == 56470 && 
b[56471] == 56471 && 
b[56472] == 56472 && 
b[56473] == 56473 && 
b[56474] == 56474 && 
b[56475] == 56475 && 
b[56476] == 56476 && 
b[56477] == 56477 && 
b[56478] == 56478 && 
b[56479] == 56479 && 
b[56480] == 56480 && 
b[56481] == 56481 && 
b[56482] == 56482 && 
b[56483] == 56483 && 
b[56484] == 56484 && 
b[56485] == 56485 && 
b[56486] == 56486 && 
b[56487] == 56487 && 
b[56488] == 56488 && 
b[56489] == 56489 && 
b[56490] == 56490 && 
b[56491] == 56491 && 
b[56492] == 56492 && 
b[56493] == 56493 && 
b[56494] == 56494 && 
b[56495] == 56495 && 
b[56496] == 56496 && 
b[56497] == 56497 && 
b[56498] == 56498 && 
b[56499] == 56499 && 
b[56500] == 56500 && 
b[56501] == 56501 && 
b[56502] == 56502 && 
b[56503] == 56503 && 
b[56504] == 56504 && 
b[56505] == 56505 && 
b[56506] == 56506 && 
b[56507] == 56507 && 
b[56508] == 56508 && 
b[56509] == 56509 && 
b[56510] == 56510 && 
b[56511] == 56511 && 
b[56512] == 56512 && 
b[56513] == 56513 && 
b[56514] == 56514 && 
b[56515] == 56515 && 
b[56516] == 56516 && 
b[56517] == 56517 && 
b[56518] == 56518 && 
b[56519] == 56519 && 
b[56520] == 56520 && 
b[56521] == 56521 && 
b[56522] == 56522 && 
b[56523] == 56523 && 
b[56524] == 56524 && 
b[56525] == 56525 && 
b[56526] == 56526 && 
b[56527] == 56527 && 
b[56528] == 56528 && 
b[56529] == 56529 && 
b[56530] == 56530 && 
b[56531] == 56531 && 
b[56532] == 56532 && 
b[56533] == 56533 && 
b[56534] == 56534 && 
b[56535] == 56535 && 
b[56536] == 56536 && 
b[56537] == 56537 && 
b[56538] == 56538 && 
b[56539] == 56539 && 
b[56540] == 56540 && 
b[56541] == 56541 && 
b[56542] == 56542 && 
b[56543] == 56543 && 
b[56544] == 56544 && 
b[56545] == 56545 && 
b[56546] == 56546 && 
b[56547] == 56547 && 
b[56548] == 56548 && 
b[56549] == 56549 && 
b[56550] == 56550 && 
b[56551] == 56551 && 
b[56552] == 56552 && 
b[56553] == 56553 && 
b[56554] == 56554 && 
b[56555] == 56555 && 
b[56556] == 56556 && 
b[56557] == 56557 && 
b[56558] == 56558 && 
b[56559] == 56559 && 
b[56560] == 56560 && 
b[56561] == 56561 && 
b[56562] == 56562 && 
b[56563] == 56563 && 
b[56564] == 56564 && 
b[56565] == 56565 && 
b[56566] == 56566 && 
b[56567] == 56567 && 
b[56568] == 56568 && 
b[56569] == 56569 && 
b[56570] == 56570 && 
b[56571] == 56571 && 
b[56572] == 56572 && 
b[56573] == 56573 && 
b[56574] == 56574 && 
b[56575] == 56575 && 
b[56576] == 56576 && 
b[56577] == 56577 && 
b[56578] == 56578 && 
b[56579] == 56579 && 
b[56580] == 56580 && 
b[56581] == 56581 && 
b[56582] == 56582 && 
b[56583] == 56583 && 
b[56584] == 56584 && 
b[56585] == 56585 && 
b[56586] == 56586 && 
b[56587] == 56587 && 
b[56588] == 56588 && 
b[56589] == 56589 && 
b[56590] == 56590 && 
b[56591] == 56591 && 
b[56592] == 56592 && 
b[56593] == 56593 && 
b[56594] == 56594 && 
b[56595] == 56595 && 
b[56596] == 56596 && 
b[56597] == 56597 && 
b[56598] == 56598 && 
b[56599] == 56599 && 
b[56600] == 56600 && 
b[56601] == 56601 && 
b[56602] == 56602 && 
b[56603] == 56603 && 
b[56604] == 56604 && 
b[56605] == 56605 && 
b[56606] == 56606 && 
b[56607] == 56607 && 
b[56608] == 56608 && 
b[56609] == 56609 && 
b[56610] == 56610 && 
b[56611] == 56611 && 
b[56612] == 56612 && 
b[56613] == 56613 && 
b[56614] == 56614 && 
b[56615] == 56615 && 
b[56616] == 56616 && 
b[56617] == 56617 && 
b[56618] == 56618 && 
b[56619] == 56619 && 
b[56620] == 56620 && 
b[56621] == 56621 && 
b[56622] == 56622 && 
b[56623] == 56623 && 
b[56624] == 56624 && 
b[56625] == 56625 && 
b[56626] == 56626 && 
b[56627] == 56627 && 
b[56628] == 56628 && 
b[56629] == 56629 && 
b[56630] == 56630 && 
b[56631] == 56631 && 
b[56632] == 56632 && 
b[56633] == 56633 && 
b[56634] == 56634 && 
b[56635] == 56635 && 
b[56636] == 56636 && 
b[56637] == 56637 && 
b[56638] == 56638 && 
b[56639] == 56639 && 
b[56640] == 56640 && 
b[56641] == 56641 && 
b[56642] == 56642 && 
b[56643] == 56643 && 
b[56644] == 56644 && 
b[56645] == 56645 && 
b[56646] == 56646 && 
b[56647] == 56647 && 
b[56648] == 56648 && 
b[56649] == 56649 && 
b[56650] == 56650 && 
b[56651] == 56651 && 
b[56652] == 56652 && 
b[56653] == 56653 && 
b[56654] == 56654 && 
b[56655] == 56655 && 
b[56656] == 56656 && 
b[56657] == 56657 && 
b[56658] == 56658 && 
b[56659] == 56659 && 
b[56660] == 56660 && 
b[56661] == 56661 && 
b[56662] == 56662 && 
b[56663] == 56663 && 
b[56664] == 56664 && 
b[56665] == 56665 && 
b[56666] == 56666 && 
b[56667] == 56667 && 
b[56668] == 56668 && 
b[56669] == 56669 && 
b[56670] == 56670 && 
b[56671] == 56671 && 
b[56672] == 56672 && 
b[56673] == 56673 && 
b[56674] == 56674 && 
b[56675] == 56675 && 
b[56676] == 56676 && 
b[56677] == 56677 && 
b[56678] == 56678 && 
b[56679] == 56679 && 
b[56680] == 56680 && 
b[56681] == 56681 && 
b[56682] == 56682 && 
b[56683] == 56683 && 
b[56684] == 56684 && 
b[56685] == 56685 && 
b[56686] == 56686 && 
b[56687] == 56687 && 
b[56688] == 56688 && 
b[56689] == 56689 && 
b[56690] == 56690 && 
b[56691] == 56691 && 
b[56692] == 56692 && 
b[56693] == 56693 && 
b[56694] == 56694 && 
b[56695] == 56695 && 
b[56696] == 56696 && 
b[56697] == 56697 && 
b[56698] == 56698 && 
b[56699] == 56699 && 
b[56700] == 56700 && 
b[56701] == 56701 && 
b[56702] == 56702 && 
b[56703] == 56703 && 
b[56704] == 56704 && 
b[56705] == 56705 && 
b[56706] == 56706 && 
b[56707] == 56707 && 
b[56708] == 56708 && 
b[56709] == 56709 && 
b[56710] == 56710 && 
b[56711] == 56711 && 
b[56712] == 56712 && 
b[56713] == 56713 && 
b[56714] == 56714 && 
b[56715] == 56715 && 
b[56716] == 56716 && 
b[56717] == 56717 && 
b[56718] == 56718 && 
b[56719] == 56719 && 
b[56720] == 56720 && 
b[56721] == 56721 && 
b[56722] == 56722 && 
b[56723] == 56723 && 
b[56724] == 56724 && 
b[56725] == 56725 && 
b[56726] == 56726 && 
b[56727] == 56727 && 
b[56728] == 56728 && 
b[56729] == 56729 && 
b[56730] == 56730 && 
b[56731] == 56731 && 
b[56732] == 56732 && 
b[56733] == 56733 && 
b[56734] == 56734 && 
b[56735] == 56735 && 
b[56736] == 56736 && 
b[56737] == 56737 && 
b[56738] == 56738 && 
b[56739] == 56739 && 
b[56740] == 56740 && 
b[56741] == 56741 && 
b[56742] == 56742 && 
b[56743] == 56743 && 
b[56744] == 56744 && 
b[56745] == 56745 && 
b[56746] == 56746 && 
b[56747] == 56747 && 
b[56748] == 56748 && 
b[56749] == 56749 && 
b[56750] == 56750 && 
b[56751] == 56751 && 
b[56752] == 56752 && 
b[56753] == 56753 && 
b[56754] == 56754 && 
b[56755] == 56755 && 
b[56756] == 56756 && 
b[56757] == 56757 && 
b[56758] == 56758 && 
b[56759] == 56759 && 
b[56760] == 56760 && 
b[56761] == 56761 && 
b[56762] == 56762 && 
b[56763] == 56763 && 
b[56764] == 56764 && 
b[56765] == 56765 && 
b[56766] == 56766 && 
b[56767] == 56767 && 
b[56768] == 56768 && 
b[56769] == 56769 && 
b[56770] == 56770 && 
b[56771] == 56771 && 
b[56772] == 56772 && 
b[56773] == 56773 && 
b[56774] == 56774 && 
b[56775] == 56775 && 
b[56776] == 56776 && 
b[56777] == 56777 && 
b[56778] == 56778 && 
b[56779] == 56779 && 
b[56780] == 56780 && 
b[56781] == 56781 && 
b[56782] == 56782 && 
b[56783] == 56783 && 
b[56784] == 56784 && 
b[56785] == 56785 && 
b[56786] == 56786 && 
b[56787] == 56787 && 
b[56788] == 56788 && 
b[56789] == 56789 && 
b[56790] == 56790 && 
b[56791] == 56791 && 
b[56792] == 56792 && 
b[56793] == 56793 && 
b[56794] == 56794 && 
b[56795] == 56795 && 
b[56796] == 56796 && 
b[56797] == 56797 && 
b[56798] == 56798 && 
b[56799] == 56799 && 
b[56800] == 56800 && 
b[56801] == 56801 && 
b[56802] == 56802 && 
b[56803] == 56803 && 
b[56804] == 56804 && 
b[56805] == 56805 && 
b[56806] == 56806 && 
b[56807] == 56807 && 
b[56808] == 56808 && 
b[56809] == 56809 && 
b[56810] == 56810 && 
b[56811] == 56811 && 
b[56812] == 56812 && 
b[56813] == 56813 && 
b[56814] == 56814 && 
b[56815] == 56815 && 
b[56816] == 56816 && 
b[56817] == 56817 && 
b[56818] == 56818 && 
b[56819] == 56819 && 
b[56820] == 56820 && 
b[56821] == 56821 && 
b[56822] == 56822 && 
b[56823] == 56823 && 
b[56824] == 56824 && 
b[56825] == 56825 && 
b[56826] == 56826 && 
b[56827] == 56827 && 
b[56828] == 56828 && 
b[56829] == 56829 && 
b[56830] == 56830 && 
b[56831] == 56831 && 
b[56832] == 56832 && 
b[56833] == 56833 && 
b[56834] == 56834 && 
b[56835] == 56835 && 
b[56836] == 56836 && 
b[56837] == 56837 && 
b[56838] == 56838 && 
b[56839] == 56839 && 
b[56840] == 56840 && 
b[56841] == 56841 && 
b[56842] == 56842 && 
b[56843] == 56843 && 
b[56844] == 56844 && 
b[56845] == 56845 && 
b[56846] == 56846 && 
b[56847] == 56847 && 
b[56848] == 56848 && 
b[56849] == 56849 && 
b[56850] == 56850 && 
b[56851] == 56851 && 
b[56852] == 56852 && 
b[56853] == 56853 && 
b[56854] == 56854 && 
b[56855] == 56855 && 
b[56856] == 56856 && 
b[56857] == 56857 && 
b[56858] == 56858 && 
b[56859] == 56859 && 
b[56860] == 56860 && 
b[56861] == 56861 && 
b[56862] == 56862 && 
b[56863] == 56863 && 
b[56864] == 56864 && 
b[56865] == 56865 && 
b[56866] == 56866 && 
b[56867] == 56867 && 
b[56868] == 56868 && 
b[56869] == 56869 && 
b[56870] == 56870 && 
b[56871] == 56871 && 
b[56872] == 56872 && 
b[56873] == 56873 && 
b[56874] == 56874 && 
b[56875] == 56875 && 
b[56876] == 56876 && 
b[56877] == 56877 && 
b[56878] == 56878 && 
b[56879] == 56879 && 
b[56880] == 56880 && 
b[56881] == 56881 && 
b[56882] == 56882 && 
b[56883] == 56883 && 
b[56884] == 56884 && 
b[56885] == 56885 && 
b[56886] == 56886 && 
b[56887] == 56887 && 
b[56888] == 56888 && 
b[56889] == 56889 && 
b[56890] == 56890 && 
b[56891] == 56891 && 
b[56892] == 56892 && 
b[56893] == 56893 && 
b[56894] == 56894 && 
b[56895] == 56895 && 
b[56896] == 56896 && 
b[56897] == 56897 && 
b[56898] == 56898 && 
b[56899] == 56899 && 
b[56900] == 56900 && 
b[56901] == 56901 && 
b[56902] == 56902 && 
b[56903] == 56903 && 
b[56904] == 56904 && 
b[56905] == 56905 && 
b[56906] == 56906 && 
b[56907] == 56907 && 
b[56908] == 56908 && 
b[56909] == 56909 && 
b[56910] == 56910 && 
b[56911] == 56911 && 
b[56912] == 56912 && 
b[56913] == 56913 && 
b[56914] == 56914 && 
b[56915] == 56915 && 
b[56916] == 56916 && 
b[56917] == 56917 && 
b[56918] == 56918 && 
b[56919] == 56919 && 
b[56920] == 56920 && 
b[56921] == 56921 && 
b[56922] == 56922 && 
b[56923] == 56923 && 
b[56924] == 56924 && 
b[56925] == 56925 && 
b[56926] == 56926 && 
b[56927] == 56927 && 
b[56928] == 56928 && 
b[56929] == 56929 && 
b[56930] == 56930 && 
b[56931] == 56931 && 
b[56932] == 56932 && 
b[56933] == 56933 && 
b[56934] == 56934 && 
b[56935] == 56935 && 
b[56936] == 56936 && 
b[56937] == 56937 && 
b[56938] == 56938 && 
b[56939] == 56939 && 
b[56940] == 56940 && 
b[56941] == 56941 && 
b[56942] == 56942 && 
b[56943] == 56943 && 
b[56944] == 56944 && 
b[56945] == 56945 && 
b[56946] == 56946 && 
b[56947] == 56947 && 
b[56948] == 56948 && 
b[56949] == 56949 && 
b[56950] == 56950 && 
b[56951] == 56951 && 
b[56952] == 56952 && 
b[56953] == 56953 && 
b[56954] == 56954 && 
b[56955] == 56955 && 
b[56956] == 56956 && 
b[56957] == 56957 && 
b[56958] == 56958 && 
b[56959] == 56959 && 
b[56960] == 56960 && 
b[56961] == 56961 && 
b[56962] == 56962 && 
b[56963] == 56963 && 
b[56964] == 56964 && 
b[56965] == 56965 && 
b[56966] == 56966 && 
b[56967] == 56967 && 
b[56968] == 56968 && 
b[56969] == 56969 && 
b[56970] == 56970 && 
b[56971] == 56971 && 
b[56972] == 56972 && 
b[56973] == 56973 && 
b[56974] == 56974 && 
b[56975] == 56975 && 
b[56976] == 56976 && 
b[56977] == 56977 && 
b[56978] == 56978 && 
b[56979] == 56979 && 
b[56980] == 56980 && 
b[56981] == 56981 && 
b[56982] == 56982 && 
b[56983] == 56983 && 
b[56984] == 56984 && 
b[56985] == 56985 && 
b[56986] == 56986 && 
b[56987] == 56987 && 
b[56988] == 56988 && 
b[56989] == 56989 && 
b[56990] == 56990 && 
b[56991] == 56991 && 
b[56992] == 56992 && 
b[56993] == 56993 && 
b[56994] == 56994 && 
b[56995] == 56995 && 
b[56996] == 56996 && 
b[56997] == 56997 && 
b[56998] == 56998 && 
b[56999] == 56999 && 
b[57000] == 57000 && 
b[57001] == 57001 && 
b[57002] == 57002 && 
b[57003] == 57003 && 
b[57004] == 57004 && 
b[57005] == 57005 && 
b[57006] == 57006 && 
b[57007] == 57007 && 
b[57008] == 57008 && 
b[57009] == 57009 && 
b[57010] == 57010 && 
b[57011] == 57011 && 
b[57012] == 57012 && 
b[57013] == 57013 && 
b[57014] == 57014 && 
b[57015] == 57015 && 
b[57016] == 57016 && 
b[57017] == 57017 && 
b[57018] == 57018 && 
b[57019] == 57019 && 
b[57020] == 57020 && 
b[57021] == 57021 && 
b[57022] == 57022 && 
b[57023] == 57023 && 
b[57024] == 57024 && 
b[57025] == 57025 && 
b[57026] == 57026 && 
b[57027] == 57027 && 
b[57028] == 57028 && 
b[57029] == 57029 && 
b[57030] == 57030 && 
b[57031] == 57031 && 
b[57032] == 57032 && 
b[57033] == 57033 && 
b[57034] == 57034 && 
b[57035] == 57035 && 
b[57036] == 57036 && 
b[57037] == 57037 && 
b[57038] == 57038 && 
b[57039] == 57039 && 
b[57040] == 57040 && 
b[57041] == 57041 && 
b[57042] == 57042 && 
b[57043] == 57043 && 
b[57044] == 57044 && 
b[57045] == 57045 && 
b[57046] == 57046 && 
b[57047] == 57047 && 
b[57048] == 57048 && 
b[57049] == 57049 && 
b[57050] == 57050 && 
b[57051] == 57051 && 
b[57052] == 57052 && 
b[57053] == 57053 && 
b[57054] == 57054 && 
b[57055] == 57055 && 
b[57056] == 57056 && 
b[57057] == 57057 && 
b[57058] == 57058 && 
b[57059] == 57059 && 
b[57060] == 57060 && 
b[57061] == 57061 && 
b[57062] == 57062 && 
b[57063] == 57063 && 
b[57064] == 57064 && 
b[57065] == 57065 && 
b[57066] == 57066 && 
b[57067] == 57067 && 
b[57068] == 57068 && 
b[57069] == 57069 && 
b[57070] == 57070 && 
b[57071] == 57071 && 
b[57072] == 57072 && 
b[57073] == 57073 && 
b[57074] == 57074 && 
b[57075] == 57075 && 
b[57076] == 57076 && 
b[57077] == 57077 && 
b[57078] == 57078 && 
b[57079] == 57079 && 
b[57080] == 57080 && 
b[57081] == 57081 && 
b[57082] == 57082 && 
b[57083] == 57083 && 
b[57084] == 57084 && 
b[57085] == 57085 && 
b[57086] == 57086 && 
b[57087] == 57087 && 
b[57088] == 57088 && 
b[57089] == 57089 && 
b[57090] == 57090 && 
b[57091] == 57091 && 
b[57092] == 57092 && 
b[57093] == 57093 && 
b[57094] == 57094 && 
b[57095] == 57095 && 
b[57096] == 57096 && 
b[57097] == 57097 && 
b[57098] == 57098 && 
b[57099] == 57099 && 
b[57100] == 57100 && 
b[57101] == 57101 && 
b[57102] == 57102 && 
b[57103] == 57103 && 
b[57104] == 57104 && 
b[57105] == 57105 && 
b[57106] == 57106 && 
b[57107] == 57107 && 
b[57108] == 57108 && 
b[57109] == 57109 && 
b[57110] == 57110 && 
b[57111] == 57111 && 
b[57112] == 57112 && 
b[57113] == 57113 && 
b[57114] == 57114 && 
b[57115] == 57115 && 
b[57116] == 57116 && 
b[57117] == 57117 && 
b[57118] == 57118 && 
b[57119] == 57119 && 
b[57120] == 57120 && 
b[57121] == 57121 && 
b[57122] == 57122 && 
b[57123] == 57123 && 
b[57124] == 57124 && 
b[57125] == 57125 && 
b[57126] == 57126 && 
b[57127] == 57127 && 
b[57128] == 57128 && 
b[57129] == 57129 && 
b[57130] == 57130 && 
b[57131] == 57131 && 
b[57132] == 57132 && 
b[57133] == 57133 && 
b[57134] == 57134 && 
b[57135] == 57135 && 
b[57136] == 57136 && 
b[57137] == 57137 && 
b[57138] == 57138 && 
b[57139] == 57139 && 
b[57140] == 57140 && 
b[57141] == 57141 && 
b[57142] == 57142 && 
b[57143] == 57143 && 
b[57144] == 57144 && 
b[57145] == 57145 && 
b[57146] == 57146 && 
b[57147] == 57147 && 
b[57148] == 57148 && 
b[57149] == 57149 && 
b[57150] == 57150 && 
b[57151] == 57151 && 
b[57152] == 57152 && 
b[57153] == 57153 && 
b[57154] == 57154 && 
b[57155] == 57155 && 
b[57156] == 57156 && 
b[57157] == 57157 && 
b[57158] == 57158 && 
b[57159] == 57159 && 
b[57160] == 57160 && 
b[57161] == 57161 && 
b[57162] == 57162 && 
b[57163] == 57163 && 
b[57164] == 57164 && 
b[57165] == 57165 && 
b[57166] == 57166 && 
b[57167] == 57167 && 
b[57168] == 57168 && 
b[57169] == 57169 && 
b[57170] == 57170 && 
b[57171] == 57171 && 
b[57172] == 57172 && 
b[57173] == 57173 && 
b[57174] == 57174 && 
b[57175] == 57175 && 
b[57176] == 57176 && 
b[57177] == 57177 && 
b[57178] == 57178 && 
b[57179] == 57179 && 
b[57180] == 57180 && 
b[57181] == 57181 && 
b[57182] == 57182 && 
b[57183] == 57183 && 
b[57184] == 57184 && 
b[57185] == 57185 && 
b[57186] == 57186 && 
b[57187] == 57187 && 
b[57188] == 57188 && 
b[57189] == 57189 && 
b[57190] == 57190 && 
b[57191] == 57191 && 
b[57192] == 57192 && 
b[57193] == 57193 && 
b[57194] == 57194 && 
b[57195] == 57195 && 
b[57196] == 57196 && 
b[57197] == 57197 && 
b[57198] == 57198 && 
b[57199] == 57199 && 
b[57200] == 57200 && 
b[57201] == 57201 && 
b[57202] == 57202 && 
b[57203] == 57203 && 
b[57204] == 57204 && 
b[57205] == 57205 && 
b[57206] == 57206 && 
b[57207] == 57207 && 
b[57208] == 57208 && 
b[57209] == 57209 && 
b[57210] == 57210 && 
b[57211] == 57211 && 
b[57212] == 57212 && 
b[57213] == 57213 && 
b[57214] == 57214 && 
b[57215] == 57215 && 
b[57216] == 57216 && 
b[57217] == 57217 && 
b[57218] == 57218 && 
b[57219] == 57219 && 
b[57220] == 57220 && 
b[57221] == 57221 && 
b[57222] == 57222 && 
b[57223] == 57223 && 
b[57224] == 57224 && 
b[57225] == 57225 && 
b[57226] == 57226 && 
b[57227] == 57227 && 
b[57228] == 57228 && 
b[57229] == 57229 && 
b[57230] == 57230 && 
b[57231] == 57231 && 
b[57232] == 57232 && 
b[57233] == 57233 && 
b[57234] == 57234 && 
b[57235] == 57235 && 
b[57236] == 57236 && 
b[57237] == 57237 && 
b[57238] == 57238 && 
b[57239] == 57239 && 
b[57240] == 57240 && 
b[57241] == 57241 && 
b[57242] == 57242 && 
b[57243] == 57243 && 
b[57244] == 57244 && 
b[57245] == 57245 && 
b[57246] == 57246 && 
b[57247] == 57247 && 
b[57248] == 57248 && 
b[57249] == 57249 && 
b[57250] == 57250 && 
b[57251] == 57251 && 
b[57252] == 57252 && 
b[57253] == 57253 && 
b[57254] == 57254 && 
b[57255] == 57255 && 
b[57256] == 57256 && 
b[57257] == 57257 && 
b[57258] == 57258 && 
b[57259] == 57259 && 
b[57260] == 57260 && 
b[57261] == 57261 && 
b[57262] == 57262 && 
b[57263] == 57263 && 
b[57264] == 57264 && 
b[57265] == 57265 && 
b[57266] == 57266 && 
b[57267] == 57267 && 
b[57268] == 57268 && 
b[57269] == 57269 && 
b[57270] == 57270 && 
b[57271] == 57271 && 
b[57272] == 57272 && 
b[57273] == 57273 && 
b[57274] == 57274 && 
b[57275] == 57275 && 
b[57276] == 57276 && 
b[57277] == 57277 && 
b[57278] == 57278 && 
b[57279] == 57279 && 
b[57280] == 57280 && 
b[57281] == 57281 && 
b[57282] == 57282 && 
b[57283] == 57283 && 
b[57284] == 57284 && 
b[57285] == 57285 && 
b[57286] == 57286 && 
b[57287] == 57287 && 
b[57288] == 57288 && 
b[57289] == 57289 && 
b[57290] == 57290 && 
b[57291] == 57291 && 
b[57292] == 57292 && 
b[57293] == 57293 && 
b[57294] == 57294 && 
b[57295] == 57295 && 
b[57296] == 57296 && 
b[57297] == 57297 && 
b[57298] == 57298 && 
b[57299] == 57299 && 
b[57300] == 57300 && 
b[57301] == 57301 && 
b[57302] == 57302 && 
b[57303] == 57303 && 
b[57304] == 57304 && 
b[57305] == 57305 && 
b[57306] == 57306 && 
b[57307] == 57307 && 
b[57308] == 57308 && 
b[57309] == 57309 && 
b[57310] == 57310 && 
b[57311] == 57311 && 
b[57312] == 57312 && 
b[57313] == 57313 && 
b[57314] == 57314 && 
b[57315] == 57315 && 
b[57316] == 57316 && 
b[57317] == 57317 && 
b[57318] == 57318 && 
b[57319] == 57319 && 
b[57320] == 57320 && 
b[57321] == 57321 && 
b[57322] == 57322 && 
b[57323] == 57323 && 
b[57324] == 57324 && 
b[57325] == 57325 && 
b[57326] == 57326 && 
b[57327] == 57327 && 
b[57328] == 57328 && 
b[57329] == 57329 && 
b[57330] == 57330 && 
b[57331] == 57331 && 
b[57332] == 57332 && 
b[57333] == 57333 && 
b[57334] == 57334 && 
b[57335] == 57335 && 
b[57336] == 57336 && 
b[57337] == 57337 && 
b[57338] == 57338 && 
b[57339] == 57339 && 
b[57340] == 57340 && 
b[57341] == 57341 && 
b[57342] == 57342 && 
b[57343] == 57343 && 
b[57344] == 57344 && 
b[57345] == 57345 && 
b[57346] == 57346 && 
b[57347] == 57347 && 
b[57348] == 57348 && 
b[57349] == 57349 && 
b[57350] == 57350 && 
b[57351] == 57351 && 
b[57352] == 57352 && 
b[57353] == 57353 && 
b[57354] == 57354 && 
b[57355] == 57355 && 
b[57356] == 57356 && 
b[57357] == 57357 && 
b[57358] == 57358 && 
b[57359] == 57359 && 
b[57360] == 57360 && 
b[57361] == 57361 && 
b[57362] == 57362 && 
b[57363] == 57363 && 
b[57364] == 57364 && 
b[57365] == 57365 && 
b[57366] == 57366 && 
b[57367] == 57367 && 
b[57368] == 57368 && 
b[57369] == 57369 && 
b[57370] == 57370 && 
b[57371] == 57371 && 
b[57372] == 57372 && 
b[57373] == 57373 && 
b[57374] == 57374 && 
b[57375] == 57375 && 
b[57376] == 57376 && 
b[57377] == 57377 && 
b[57378] == 57378 && 
b[57379] == 57379 && 
b[57380] == 57380 && 
b[57381] == 57381 && 
b[57382] == 57382 && 
b[57383] == 57383 && 
b[57384] == 57384 && 
b[57385] == 57385 && 
b[57386] == 57386 && 
b[57387] == 57387 && 
b[57388] == 57388 && 
b[57389] == 57389 && 
b[57390] == 57390 && 
b[57391] == 57391 && 
b[57392] == 57392 && 
b[57393] == 57393 && 
b[57394] == 57394 && 
b[57395] == 57395 && 
b[57396] == 57396 && 
b[57397] == 57397 && 
b[57398] == 57398 && 
b[57399] == 57399 && 
b[57400] == 57400 && 
b[57401] == 57401 && 
b[57402] == 57402 && 
b[57403] == 57403 && 
b[57404] == 57404 && 
b[57405] == 57405 && 
b[57406] == 57406 && 
b[57407] == 57407 && 
b[57408] == 57408 && 
b[57409] == 57409 && 
b[57410] == 57410 && 
b[57411] == 57411 && 
b[57412] == 57412 && 
b[57413] == 57413 && 
b[57414] == 57414 && 
b[57415] == 57415 && 
b[57416] == 57416 && 
b[57417] == 57417 && 
b[57418] == 57418 && 
b[57419] == 57419 && 
b[57420] == 57420 && 
b[57421] == 57421 && 
b[57422] == 57422 && 
b[57423] == 57423 && 
b[57424] == 57424 && 
b[57425] == 57425 && 
b[57426] == 57426 && 
b[57427] == 57427 && 
b[57428] == 57428 && 
b[57429] == 57429 && 
b[57430] == 57430 && 
b[57431] == 57431 && 
b[57432] == 57432 && 
b[57433] == 57433 && 
b[57434] == 57434 && 
b[57435] == 57435 && 
b[57436] == 57436 && 
b[57437] == 57437 && 
b[57438] == 57438 && 
b[57439] == 57439 && 
b[57440] == 57440 && 
b[57441] == 57441 && 
b[57442] == 57442 && 
b[57443] == 57443 && 
b[57444] == 57444 && 
b[57445] == 57445 && 
b[57446] == 57446 && 
b[57447] == 57447 && 
b[57448] == 57448 && 
b[57449] == 57449 && 
b[57450] == 57450 && 
b[57451] == 57451 && 
b[57452] == 57452 && 
b[57453] == 57453 && 
b[57454] == 57454 && 
b[57455] == 57455 && 
b[57456] == 57456 && 
b[57457] == 57457 && 
b[57458] == 57458 && 
b[57459] == 57459 && 
b[57460] == 57460 && 
b[57461] == 57461 && 
b[57462] == 57462 && 
b[57463] == 57463 && 
b[57464] == 57464 && 
b[57465] == 57465 && 
b[57466] == 57466 && 
b[57467] == 57467 && 
b[57468] == 57468 && 
b[57469] == 57469 && 
b[57470] == 57470 && 
b[57471] == 57471 && 
b[57472] == 57472 && 
b[57473] == 57473 && 
b[57474] == 57474 && 
b[57475] == 57475 && 
b[57476] == 57476 && 
b[57477] == 57477 && 
b[57478] == 57478 && 
b[57479] == 57479 && 
b[57480] == 57480 && 
b[57481] == 57481 && 
b[57482] == 57482 && 
b[57483] == 57483 && 
b[57484] == 57484 && 
b[57485] == 57485 && 
b[57486] == 57486 && 
b[57487] == 57487 && 
b[57488] == 57488 && 
b[57489] == 57489 && 
b[57490] == 57490 && 
b[57491] == 57491 && 
b[57492] == 57492 && 
b[57493] == 57493 && 
b[57494] == 57494 && 
b[57495] == 57495 && 
b[57496] == 57496 && 
b[57497] == 57497 && 
b[57498] == 57498 && 
b[57499] == 57499 && 
b[57500] == 57500 && 
b[57501] == 57501 && 
b[57502] == 57502 && 
b[57503] == 57503 && 
b[57504] == 57504 && 
b[57505] == 57505 && 
b[57506] == 57506 && 
b[57507] == 57507 && 
b[57508] == 57508 && 
b[57509] == 57509 && 
b[57510] == 57510 && 
b[57511] == 57511 && 
b[57512] == 57512 && 
b[57513] == 57513 && 
b[57514] == 57514 && 
b[57515] == 57515 && 
b[57516] == 57516 && 
b[57517] == 57517 && 
b[57518] == 57518 && 
b[57519] == 57519 && 
b[57520] == 57520 && 
b[57521] == 57521 && 
b[57522] == 57522 && 
b[57523] == 57523 && 
b[57524] == 57524 && 
b[57525] == 57525 && 
b[57526] == 57526 && 
b[57527] == 57527 && 
b[57528] == 57528 && 
b[57529] == 57529 && 
b[57530] == 57530 && 
b[57531] == 57531 && 
b[57532] == 57532 && 
b[57533] == 57533 && 
b[57534] == 57534 && 
b[57535] == 57535 && 
b[57536] == 57536 && 
b[57537] == 57537 && 
b[57538] == 57538 && 
b[57539] == 57539 && 
b[57540] == 57540 && 
b[57541] == 57541 && 
b[57542] == 57542 && 
b[57543] == 57543 && 
b[57544] == 57544 && 
b[57545] == 57545 && 
b[57546] == 57546 && 
b[57547] == 57547 && 
b[57548] == 57548 && 
b[57549] == 57549 && 
b[57550] == 57550 && 
b[57551] == 57551 && 
b[57552] == 57552 && 
b[57553] == 57553 && 
b[57554] == 57554 && 
b[57555] == 57555 && 
b[57556] == 57556 && 
b[57557] == 57557 && 
b[57558] == 57558 && 
b[57559] == 57559 && 
b[57560] == 57560 && 
b[57561] == 57561 && 
b[57562] == 57562 && 
b[57563] == 57563 && 
b[57564] == 57564 && 
b[57565] == 57565 && 
b[57566] == 57566 && 
b[57567] == 57567 && 
b[57568] == 57568 && 
b[57569] == 57569 && 
b[57570] == 57570 && 
b[57571] == 57571 && 
b[57572] == 57572 && 
b[57573] == 57573 && 
b[57574] == 57574 && 
b[57575] == 57575 && 
b[57576] == 57576 && 
b[57577] == 57577 && 
b[57578] == 57578 && 
b[57579] == 57579 && 
b[57580] == 57580 && 
b[57581] == 57581 && 
b[57582] == 57582 && 
b[57583] == 57583 && 
b[57584] == 57584 && 
b[57585] == 57585 && 
b[57586] == 57586 && 
b[57587] == 57587 && 
b[57588] == 57588 && 
b[57589] == 57589 && 
b[57590] == 57590 && 
b[57591] == 57591 && 
b[57592] == 57592 && 
b[57593] == 57593 && 
b[57594] == 57594 && 
b[57595] == 57595 && 
b[57596] == 57596 && 
b[57597] == 57597 && 
b[57598] == 57598 && 
b[57599] == 57599 && 
b[57600] == 57600 && 
b[57601] == 57601 && 
b[57602] == 57602 && 
b[57603] == 57603 && 
b[57604] == 57604 && 
b[57605] == 57605 && 
b[57606] == 57606 && 
b[57607] == 57607 && 
b[57608] == 57608 && 
b[57609] == 57609 && 
b[57610] == 57610 && 
b[57611] == 57611 && 
b[57612] == 57612 && 
b[57613] == 57613 && 
b[57614] == 57614 && 
b[57615] == 57615 && 
b[57616] == 57616 && 
b[57617] == 57617 && 
b[57618] == 57618 && 
b[57619] == 57619 && 
b[57620] == 57620 && 
b[57621] == 57621 && 
b[57622] == 57622 && 
b[57623] == 57623 && 
b[57624] == 57624 && 
b[57625] == 57625 && 
b[57626] == 57626 && 
b[57627] == 57627 && 
b[57628] == 57628 && 
b[57629] == 57629 && 
b[57630] == 57630 && 
b[57631] == 57631 && 
b[57632] == 57632 && 
b[57633] == 57633 && 
b[57634] == 57634 && 
b[57635] == 57635 && 
b[57636] == 57636 && 
b[57637] == 57637 && 
b[57638] == 57638 && 
b[57639] == 57639 && 
b[57640] == 57640 && 
b[57641] == 57641 && 
b[57642] == 57642 && 
b[57643] == 57643 && 
b[57644] == 57644 && 
b[57645] == 57645 && 
b[57646] == 57646 && 
b[57647] == 57647 && 
b[57648] == 57648 && 
b[57649] == 57649 && 
b[57650] == 57650 && 
b[57651] == 57651 && 
b[57652] == 57652 && 
b[57653] == 57653 && 
b[57654] == 57654 && 
b[57655] == 57655 && 
b[57656] == 57656 && 
b[57657] == 57657 && 
b[57658] == 57658 && 
b[57659] == 57659 && 
b[57660] == 57660 && 
b[57661] == 57661 && 
b[57662] == 57662 && 
b[57663] == 57663 && 
b[57664] == 57664 && 
b[57665] == 57665 && 
b[57666] == 57666 && 
b[57667] == 57667 && 
b[57668] == 57668 && 
b[57669] == 57669 && 
b[57670] == 57670 && 
b[57671] == 57671 && 
b[57672] == 57672 && 
b[57673] == 57673 && 
b[57674] == 57674 && 
b[57675] == 57675 && 
b[57676] == 57676 && 
b[57677] == 57677 && 
b[57678] == 57678 && 
b[57679] == 57679 && 
b[57680] == 57680 && 
b[57681] == 57681 && 
b[57682] == 57682 && 
b[57683] == 57683 && 
b[57684] == 57684 && 
b[57685] == 57685 && 
b[57686] == 57686 && 
b[57687] == 57687 && 
b[57688] == 57688 && 
b[57689] == 57689 && 
b[57690] == 57690 && 
b[57691] == 57691 && 
b[57692] == 57692 && 
b[57693] == 57693 && 
b[57694] == 57694 && 
b[57695] == 57695 && 
b[57696] == 57696 && 
b[57697] == 57697 && 
b[57698] == 57698 && 
b[57699] == 57699 && 
b[57700] == 57700 && 
b[57701] == 57701 && 
b[57702] == 57702 && 
b[57703] == 57703 && 
b[57704] == 57704 && 
b[57705] == 57705 && 
b[57706] == 57706 && 
b[57707] == 57707 && 
b[57708] == 57708 && 
b[57709] == 57709 && 
b[57710] == 57710 && 
b[57711] == 57711 && 
b[57712] == 57712 && 
b[57713] == 57713 && 
b[57714] == 57714 && 
b[57715] == 57715 && 
b[57716] == 57716 && 
b[57717] == 57717 && 
b[57718] == 57718 && 
b[57719] == 57719 && 
b[57720] == 57720 && 
b[57721] == 57721 && 
b[57722] == 57722 && 
b[57723] == 57723 && 
b[57724] == 57724 && 
b[57725] == 57725 && 
b[57726] == 57726 && 
b[57727] == 57727 && 
b[57728] == 57728 && 
b[57729] == 57729 && 
b[57730] == 57730 && 
b[57731] == 57731 && 
b[57732] == 57732 && 
b[57733] == 57733 && 
b[57734] == 57734 && 
b[57735] == 57735 && 
b[57736] == 57736 && 
b[57737] == 57737 && 
b[57738] == 57738 && 
b[57739] == 57739 && 
b[57740] == 57740 && 
b[57741] == 57741 && 
b[57742] == 57742 && 
b[57743] == 57743 && 
b[57744] == 57744 && 
b[57745] == 57745 && 
b[57746] == 57746 && 
b[57747] == 57747 && 
b[57748] == 57748 && 
b[57749] == 57749 && 
b[57750] == 57750 && 
b[57751] == 57751 && 
b[57752] == 57752 && 
b[57753] == 57753 && 
b[57754] == 57754 && 
b[57755] == 57755 && 
b[57756] == 57756 && 
b[57757] == 57757 && 
b[57758] == 57758 && 
b[57759] == 57759 && 
b[57760] == 57760 && 
b[57761] == 57761 && 
b[57762] == 57762 && 
b[57763] == 57763 && 
b[57764] == 57764 && 
b[57765] == 57765 && 
b[57766] == 57766 && 
b[57767] == 57767 && 
b[57768] == 57768 && 
b[57769] == 57769 && 
b[57770] == 57770 && 
b[57771] == 57771 && 
b[57772] == 57772 && 
b[57773] == 57773 && 
b[57774] == 57774 && 
b[57775] == 57775 && 
b[57776] == 57776 && 
b[57777] == 57777 && 
b[57778] == 57778 && 
b[57779] == 57779 && 
b[57780] == 57780 && 
b[57781] == 57781 && 
b[57782] == 57782 && 
b[57783] == 57783 && 
b[57784] == 57784 && 
b[57785] == 57785 && 
b[57786] == 57786 && 
b[57787] == 57787 && 
b[57788] == 57788 && 
b[57789] == 57789 && 
b[57790] == 57790 && 
b[57791] == 57791 && 
b[57792] == 57792 && 
b[57793] == 57793 && 
b[57794] == 57794 && 
b[57795] == 57795 && 
b[57796] == 57796 && 
b[57797] == 57797 && 
b[57798] == 57798 && 
b[57799] == 57799 && 
b[57800] == 57800 && 
b[57801] == 57801 && 
b[57802] == 57802 && 
b[57803] == 57803 && 
b[57804] == 57804 && 
b[57805] == 57805 && 
b[57806] == 57806 && 
b[57807] == 57807 && 
b[57808] == 57808 && 
b[57809] == 57809 && 
b[57810] == 57810 && 
b[57811] == 57811 && 
b[57812] == 57812 && 
b[57813] == 57813 && 
b[57814] == 57814 && 
b[57815] == 57815 && 
b[57816] == 57816 && 
b[57817] == 57817 && 
b[57818] == 57818 && 
b[57819] == 57819 && 
b[57820] == 57820 && 
b[57821] == 57821 && 
b[57822] == 57822 && 
b[57823] == 57823 && 
b[57824] == 57824 && 
b[57825] == 57825 && 
b[57826] == 57826 && 
b[57827] == 57827 && 
b[57828] == 57828 && 
b[57829] == 57829 && 
b[57830] == 57830 && 
b[57831] == 57831 && 
b[57832] == 57832 && 
b[57833] == 57833 && 
b[57834] == 57834 && 
b[57835] == 57835 && 
b[57836] == 57836 && 
b[57837] == 57837 && 
b[57838] == 57838 && 
b[57839] == 57839 && 
b[57840] == 57840 && 
b[57841] == 57841 && 
b[57842] == 57842 && 
b[57843] == 57843 && 
b[57844] == 57844 && 
b[57845] == 57845 && 
b[57846] == 57846 && 
b[57847] == 57847 && 
b[57848] == 57848 && 
b[57849] == 57849 && 
b[57850] == 57850 && 
b[57851] == 57851 && 
b[57852] == 57852 && 
b[57853] == 57853 && 
b[57854] == 57854 && 
b[57855] == 57855 && 
b[57856] == 57856 && 
b[57857] == 57857 && 
b[57858] == 57858 && 
b[57859] == 57859 && 
b[57860] == 57860 && 
b[57861] == 57861 && 
b[57862] == 57862 && 
b[57863] == 57863 && 
b[57864] == 57864 && 
b[57865] == 57865 && 
b[57866] == 57866 && 
b[57867] == 57867 && 
b[57868] == 57868 && 
b[57869] == 57869 && 
b[57870] == 57870 && 
b[57871] == 57871 && 
b[57872] == 57872 && 
b[57873] == 57873 && 
b[57874] == 57874 && 
b[57875] == 57875 && 
b[57876] == 57876 && 
b[57877] == 57877 && 
b[57878] == 57878 && 
b[57879] == 57879 && 
b[57880] == 57880 && 
b[57881] == 57881 && 
b[57882] == 57882 && 
b[57883] == 57883 && 
b[57884] == 57884 && 
b[57885] == 57885 && 
b[57886] == 57886 && 
b[57887] == 57887 && 
b[57888] == 57888 && 
b[57889] == 57889 && 
b[57890] == 57890 && 
b[57891] == 57891 && 
b[57892] == 57892 && 
b[57893] == 57893 && 
b[57894] == 57894 && 
b[57895] == 57895 && 
b[57896] == 57896 && 
b[57897] == 57897 && 
b[57898] == 57898 && 
b[57899] == 57899 && 
b[57900] == 57900 && 
b[57901] == 57901 && 
b[57902] == 57902 && 
b[57903] == 57903 && 
b[57904] == 57904 && 
b[57905] == 57905 && 
b[57906] == 57906 && 
b[57907] == 57907 && 
b[57908] == 57908 && 
b[57909] == 57909 && 
b[57910] == 57910 && 
b[57911] == 57911 && 
b[57912] == 57912 && 
b[57913] == 57913 && 
b[57914] == 57914 && 
b[57915] == 57915 && 
b[57916] == 57916 && 
b[57917] == 57917 && 
b[57918] == 57918 && 
b[57919] == 57919 && 
b[57920] == 57920 && 
b[57921] == 57921 && 
b[57922] == 57922 && 
b[57923] == 57923 && 
b[57924] == 57924 && 
b[57925] == 57925 && 
b[57926] == 57926 && 
b[57927] == 57927 && 
b[57928] == 57928 && 
b[57929] == 57929 && 
b[57930] == 57930 && 
b[57931] == 57931 && 
b[57932] == 57932 && 
b[57933] == 57933 && 
b[57934] == 57934 && 
b[57935] == 57935 && 
b[57936] == 57936 && 
b[57937] == 57937 && 
b[57938] == 57938 && 
b[57939] == 57939 && 
b[57940] == 57940 && 
b[57941] == 57941 && 
b[57942] == 57942 && 
b[57943] == 57943 && 
b[57944] == 57944 && 
b[57945] == 57945 && 
b[57946] == 57946 && 
b[57947] == 57947 && 
b[57948] == 57948 && 
b[57949] == 57949 && 
b[57950] == 57950 && 
b[57951] == 57951 && 
b[57952] == 57952 && 
b[57953] == 57953 && 
b[57954] == 57954 && 
b[57955] == 57955 && 
b[57956] == 57956 && 
b[57957] == 57957 && 
b[57958] == 57958 && 
b[57959] == 57959 && 
b[57960] == 57960 && 
b[57961] == 57961 && 
b[57962] == 57962 && 
b[57963] == 57963 && 
b[57964] == 57964 && 
b[57965] == 57965 && 
b[57966] == 57966 && 
b[57967] == 57967 && 
b[57968] == 57968 && 
b[57969] == 57969 && 
b[57970] == 57970 && 
b[57971] == 57971 && 
b[57972] == 57972 && 
b[57973] == 57973 && 
b[57974] == 57974 && 
b[57975] == 57975 && 
b[57976] == 57976 && 
b[57977] == 57977 && 
b[57978] == 57978 && 
b[57979] == 57979 && 
b[57980] == 57980 && 
b[57981] == 57981 && 
b[57982] == 57982 && 
b[57983] == 57983 && 
b[57984] == 57984 && 
b[57985] == 57985 && 
b[57986] == 57986 && 
b[57987] == 57987 && 
b[57988] == 57988 && 
b[57989] == 57989 && 
b[57990] == 57990 && 
b[57991] == 57991 && 
b[57992] == 57992 && 
b[57993] == 57993 && 
b[57994] == 57994 && 
b[57995] == 57995 && 
b[57996] == 57996 && 
b[57997] == 57997 && 
b[57998] == 57998 && 
b[57999] == 57999 && 
b[58000] == 58000 && 
b[58001] == 58001 && 
b[58002] == 58002 && 
b[58003] == 58003 && 
b[58004] == 58004 && 
b[58005] == 58005 && 
b[58006] == 58006 && 
b[58007] == 58007 && 
b[58008] == 58008 && 
b[58009] == 58009 && 
b[58010] == 58010 && 
b[58011] == 58011 && 
b[58012] == 58012 && 
b[58013] == 58013 && 
b[58014] == 58014 && 
b[58015] == 58015 && 
b[58016] == 58016 && 
b[58017] == 58017 && 
b[58018] == 58018 && 
b[58019] == 58019 && 
b[58020] == 58020 && 
b[58021] == 58021 && 
b[58022] == 58022 && 
b[58023] == 58023 && 
b[58024] == 58024 && 
b[58025] == 58025 && 
b[58026] == 58026 && 
b[58027] == 58027 && 
b[58028] == 58028 && 
b[58029] == 58029 && 
b[58030] == 58030 && 
b[58031] == 58031 && 
b[58032] == 58032 && 
b[58033] == 58033 && 
b[58034] == 58034 && 
b[58035] == 58035 && 
b[58036] == 58036 && 
b[58037] == 58037 && 
b[58038] == 58038 && 
b[58039] == 58039 && 
b[58040] == 58040 && 
b[58041] == 58041 && 
b[58042] == 58042 && 
b[58043] == 58043 && 
b[58044] == 58044 && 
b[58045] == 58045 && 
b[58046] == 58046 && 
b[58047] == 58047 && 
b[58048] == 58048 && 
b[58049] == 58049 && 
b[58050] == 58050 && 
b[58051] == 58051 && 
b[58052] == 58052 && 
b[58053] == 58053 && 
b[58054] == 58054 && 
b[58055] == 58055 && 
b[58056] == 58056 && 
b[58057] == 58057 && 
b[58058] == 58058 && 
b[58059] == 58059 && 
b[58060] == 58060 && 
b[58061] == 58061 && 
b[58062] == 58062 && 
b[58063] == 58063 && 
b[58064] == 58064 && 
b[58065] == 58065 && 
b[58066] == 58066 && 
b[58067] == 58067 && 
b[58068] == 58068 && 
b[58069] == 58069 && 
b[58070] == 58070 && 
b[58071] == 58071 && 
b[58072] == 58072 && 
b[58073] == 58073 && 
b[58074] == 58074 && 
b[58075] == 58075 && 
b[58076] == 58076 && 
b[58077] == 58077 && 
b[58078] == 58078 && 
b[58079] == 58079 && 
b[58080] == 58080 && 
b[58081] == 58081 && 
b[58082] == 58082 && 
b[58083] == 58083 && 
b[58084] == 58084 && 
b[58085] == 58085 && 
b[58086] == 58086 && 
b[58087] == 58087 && 
b[58088] == 58088 && 
b[58089] == 58089 && 
b[58090] == 58090 && 
b[58091] == 58091 && 
b[58092] == 58092 && 
b[58093] == 58093 && 
b[58094] == 58094 && 
b[58095] == 58095 && 
b[58096] == 58096 && 
b[58097] == 58097 && 
b[58098] == 58098 && 
b[58099] == 58099 && 
b[58100] == 58100 && 
b[58101] == 58101 && 
b[58102] == 58102 && 
b[58103] == 58103 && 
b[58104] == 58104 && 
b[58105] == 58105 && 
b[58106] == 58106 && 
b[58107] == 58107 && 
b[58108] == 58108 && 
b[58109] == 58109 && 
b[58110] == 58110 && 
b[58111] == 58111 && 
b[58112] == 58112 && 
b[58113] == 58113 && 
b[58114] == 58114 && 
b[58115] == 58115 && 
b[58116] == 58116 && 
b[58117] == 58117 && 
b[58118] == 58118 && 
b[58119] == 58119 && 
b[58120] == 58120 && 
b[58121] == 58121 && 
b[58122] == 58122 && 
b[58123] == 58123 && 
b[58124] == 58124 && 
b[58125] == 58125 && 
b[58126] == 58126 && 
b[58127] == 58127 && 
b[58128] == 58128 && 
b[58129] == 58129 && 
b[58130] == 58130 && 
b[58131] == 58131 && 
b[58132] == 58132 && 
b[58133] == 58133 && 
b[58134] == 58134 && 
b[58135] == 58135 && 
b[58136] == 58136 && 
b[58137] == 58137 && 
b[58138] == 58138 && 
b[58139] == 58139 && 
b[58140] == 58140 && 
b[58141] == 58141 && 
b[58142] == 58142 && 
b[58143] == 58143 && 
b[58144] == 58144 && 
b[58145] == 58145 && 
b[58146] == 58146 && 
b[58147] == 58147 && 
b[58148] == 58148 && 
b[58149] == 58149 && 
b[58150] == 58150 && 
b[58151] == 58151 && 
b[58152] == 58152 && 
b[58153] == 58153 && 
b[58154] == 58154 && 
b[58155] == 58155 && 
b[58156] == 58156 && 
b[58157] == 58157 && 
b[58158] == 58158 && 
b[58159] == 58159 && 
b[58160] == 58160 && 
b[58161] == 58161 && 
b[58162] == 58162 && 
b[58163] == 58163 && 
b[58164] == 58164 && 
b[58165] == 58165 && 
b[58166] == 58166 && 
b[58167] == 58167 && 
b[58168] == 58168 && 
b[58169] == 58169 && 
b[58170] == 58170 && 
b[58171] == 58171 && 
b[58172] == 58172 && 
b[58173] == 58173 && 
b[58174] == 58174 && 
b[58175] == 58175 && 
b[58176] == 58176 && 
b[58177] == 58177 && 
b[58178] == 58178 && 
b[58179] == 58179 && 
b[58180] == 58180 && 
b[58181] == 58181 && 
b[58182] == 58182 && 
b[58183] == 58183 && 
b[58184] == 58184 && 
b[58185] == 58185 && 
b[58186] == 58186 && 
b[58187] == 58187 && 
b[58188] == 58188 && 
b[58189] == 58189 && 
b[58190] == 58190 && 
b[58191] == 58191 && 
b[58192] == 58192 && 
b[58193] == 58193 && 
b[58194] == 58194 && 
b[58195] == 58195 && 
b[58196] == 58196 && 
b[58197] == 58197 && 
b[58198] == 58198 && 
b[58199] == 58199 && 
b[58200] == 58200 && 
b[58201] == 58201 && 
b[58202] == 58202 && 
b[58203] == 58203 && 
b[58204] == 58204 && 
b[58205] == 58205 && 
b[58206] == 58206 && 
b[58207] == 58207 && 
b[58208] == 58208 && 
b[58209] == 58209 && 
b[58210] == 58210 && 
b[58211] == 58211 && 
b[58212] == 58212 && 
b[58213] == 58213 && 
b[58214] == 58214 && 
b[58215] == 58215 && 
b[58216] == 58216 && 
b[58217] == 58217 && 
b[58218] == 58218 && 
b[58219] == 58219 && 
b[58220] == 58220 && 
b[58221] == 58221 && 
b[58222] == 58222 && 
b[58223] == 58223 && 
b[58224] == 58224 && 
b[58225] == 58225 && 
b[58226] == 58226 && 
b[58227] == 58227 && 
b[58228] == 58228 && 
b[58229] == 58229 && 
b[58230] == 58230 && 
b[58231] == 58231 && 
b[58232] == 58232 && 
b[58233] == 58233 && 
b[58234] == 58234 && 
b[58235] == 58235 && 
b[58236] == 58236 && 
b[58237] == 58237 && 
b[58238] == 58238 && 
b[58239] == 58239 && 
b[58240] == 58240 && 
b[58241] == 58241 && 
b[58242] == 58242 && 
b[58243] == 58243 && 
b[58244] == 58244 && 
b[58245] == 58245 && 
b[58246] == 58246 && 
b[58247] == 58247 && 
b[58248] == 58248 && 
b[58249] == 58249 && 
b[58250] == 58250 && 
b[58251] == 58251 && 
b[58252] == 58252 && 
b[58253] == 58253 && 
b[58254] == 58254 && 
b[58255] == 58255 && 
b[58256] == 58256 && 
b[58257] == 58257 && 
b[58258] == 58258 && 
b[58259] == 58259 && 
b[58260] == 58260 && 
b[58261] == 58261 && 
b[58262] == 58262 && 
b[58263] == 58263 && 
b[58264] == 58264 && 
b[58265] == 58265 && 
b[58266] == 58266 && 
b[58267] == 58267 && 
b[58268] == 58268 && 
b[58269] == 58269 && 
b[58270] == 58270 && 
b[58271] == 58271 && 
b[58272] == 58272 && 
b[58273] == 58273 && 
b[58274] == 58274 && 
b[58275] == 58275 && 
b[58276] == 58276 && 
b[58277] == 58277 && 
b[58278] == 58278 && 
b[58279] == 58279 && 
b[58280] == 58280 && 
b[58281] == 58281 && 
b[58282] == 58282 && 
b[58283] == 58283 && 
b[58284] == 58284 && 
b[58285] == 58285 && 
b[58286] == 58286 && 
b[58287] == 58287 && 
b[58288] == 58288 && 
b[58289] == 58289 && 
b[58290] == 58290 && 
b[58291] == 58291 && 
b[58292] == 58292 && 
b[58293] == 58293 && 
b[58294] == 58294 && 
b[58295] == 58295 && 
b[58296] == 58296 && 
b[58297] == 58297 && 
b[58298] == 58298 && 
b[58299] == 58299 && 
b[58300] == 58300 && 
b[58301] == 58301 && 
b[58302] == 58302 && 
b[58303] == 58303 && 
b[58304] == 58304 && 
b[58305] == 58305 && 
b[58306] == 58306 && 
b[58307] == 58307 && 
b[58308] == 58308 && 
b[58309] == 58309 && 
b[58310] == 58310 && 
b[58311] == 58311 && 
b[58312] == 58312 && 
b[58313] == 58313 && 
b[58314] == 58314 && 
b[58315] == 58315 && 
b[58316] == 58316 && 
b[58317] == 58317 && 
b[58318] == 58318 && 
b[58319] == 58319 && 
b[58320] == 58320 && 
b[58321] == 58321 && 
b[58322] == 58322 && 
b[58323] == 58323 && 
b[58324] == 58324 && 
b[58325] == 58325 && 
b[58326] == 58326 && 
b[58327] == 58327 && 
b[58328] == 58328 && 
b[58329] == 58329 && 
b[58330] == 58330 && 
b[58331] == 58331 && 
b[58332] == 58332 && 
b[58333] == 58333 && 
b[58334] == 58334 && 
b[58335] == 58335 && 
b[58336] == 58336 && 
b[58337] == 58337 && 
b[58338] == 58338 && 
b[58339] == 58339 && 
b[58340] == 58340 && 
b[58341] == 58341 && 
b[58342] == 58342 && 
b[58343] == 58343 && 
b[58344] == 58344 && 
b[58345] == 58345 && 
b[58346] == 58346 && 
b[58347] == 58347 && 
b[58348] == 58348 && 
b[58349] == 58349 && 
b[58350] == 58350 && 
b[58351] == 58351 && 
b[58352] == 58352 && 
b[58353] == 58353 && 
b[58354] == 58354 && 
b[58355] == 58355 && 
b[58356] == 58356 && 
b[58357] == 58357 && 
b[58358] == 58358 && 
b[58359] == 58359 && 
b[58360] == 58360 && 
b[58361] == 58361 && 
b[58362] == 58362 && 
b[58363] == 58363 && 
b[58364] == 58364 && 
b[58365] == 58365 && 
b[58366] == 58366 && 
b[58367] == 58367 && 
b[58368] == 58368 && 
b[58369] == 58369 && 
b[58370] == 58370 && 
b[58371] == 58371 && 
b[58372] == 58372 && 
b[58373] == 58373 && 
b[58374] == 58374 && 
b[58375] == 58375 && 
b[58376] == 58376 && 
b[58377] == 58377 && 
b[58378] == 58378 && 
b[58379] == 58379 && 
b[58380] == 58380 && 
b[58381] == 58381 && 
b[58382] == 58382 && 
b[58383] == 58383 && 
b[58384] == 58384 && 
b[58385] == 58385 && 
b[58386] == 58386 && 
b[58387] == 58387 && 
b[58388] == 58388 && 
b[58389] == 58389 && 
b[58390] == 58390 && 
b[58391] == 58391 && 
b[58392] == 58392 && 
b[58393] == 58393 && 
b[58394] == 58394 && 
b[58395] == 58395 && 
b[58396] == 58396 && 
b[58397] == 58397 && 
b[58398] == 58398 && 
b[58399] == 58399 && 
b[58400] == 58400 && 
b[58401] == 58401 && 
b[58402] == 58402 && 
b[58403] == 58403 && 
b[58404] == 58404 && 
b[58405] == 58405 && 
b[58406] == 58406 && 
b[58407] == 58407 && 
b[58408] == 58408 && 
b[58409] == 58409 && 
b[58410] == 58410 && 
b[58411] == 58411 && 
b[58412] == 58412 && 
b[58413] == 58413 && 
b[58414] == 58414 && 
b[58415] == 58415 && 
b[58416] == 58416 && 
b[58417] == 58417 && 
b[58418] == 58418 && 
b[58419] == 58419 && 
b[58420] == 58420 && 
b[58421] == 58421 && 
b[58422] == 58422 && 
b[58423] == 58423 && 
b[58424] == 58424 && 
b[58425] == 58425 && 
b[58426] == 58426 && 
b[58427] == 58427 && 
b[58428] == 58428 && 
b[58429] == 58429 && 
b[58430] == 58430 && 
b[58431] == 58431 && 
b[58432] == 58432 && 
b[58433] == 58433 && 
b[58434] == 58434 && 
b[58435] == 58435 && 
b[58436] == 58436 && 
b[58437] == 58437 && 
b[58438] == 58438 && 
b[58439] == 58439 && 
b[58440] == 58440 && 
b[58441] == 58441 && 
b[58442] == 58442 && 
b[58443] == 58443 && 
b[58444] == 58444 && 
b[58445] == 58445 && 
b[58446] == 58446 && 
b[58447] == 58447 && 
b[58448] == 58448 && 
b[58449] == 58449 && 
b[58450] == 58450 && 
b[58451] == 58451 && 
b[58452] == 58452 && 
b[58453] == 58453 && 
b[58454] == 58454 && 
b[58455] == 58455 && 
b[58456] == 58456 && 
b[58457] == 58457 && 
b[58458] == 58458 && 
b[58459] == 58459 && 
b[58460] == 58460 && 
b[58461] == 58461 && 
b[58462] == 58462 && 
b[58463] == 58463 && 
b[58464] == 58464 && 
b[58465] == 58465 && 
b[58466] == 58466 && 
b[58467] == 58467 && 
b[58468] == 58468 && 
b[58469] == 58469 && 
b[58470] == 58470 && 
b[58471] == 58471 && 
b[58472] == 58472 && 
b[58473] == 58473 && 
b[58474] == 58474 && 
b[58475] == 58475 && 
b[58476] == 58476 && 
b[58477] == 58477 && 
b[58478] == 58478 && 
b[58479] == 58479 && 
b[58480] == 58480 && 
b[58481] == 58481 && 
b[58482] == 58482 && 
b[58483] == 58483 && 
b[58484] == 58484 && 
b[58485] == 58485 && 
b[58486] == 58486 && 
b[58487] == 58487 && 
b[58488] == 58488 && 
b[58489] == 58489 && 
b[58490] == 58490 && 
b[58491] == 58491 && 
b[58492] == 58492 && 
b[58493] == 58493 && 
b[58494] == 58494 && 
b[58495] == 58495 && 
b[58496] == 58496 && 
b[58497] == 58497 && 
b[58498] == 58498 && 
b[58499] == 58499 && 
b[58500] == 58500 && 
b[58501] == 58501 && 
b[58502] == 58502 && 
b[58503] == 58503 && 
b[58504] == 58504 && 
b[58505] == 58505 && 
b[58506] == 58506 && 
b[58507] == 58507 && 
b[58508] == 58508 && 
b[58509] == 58509 && 
b[58510] == 58510 && 
b[58511] == 58511 && 
b[58512] == 58512 && 
b[58513] == 58513 && 
b[58514] == 58514 && 
b[58515] == 58515 && 
b[58516] == 58516 && 
b[58517] == 58517 && 
b[58518] == 58518 && 
b[58519] == 58519 && 
b[58520] == 58520 && 
b[58521] == 58521 && 
b[58522] == 58522 && 
b[58523] == 58523 && 
b[58524] == 58524 && 
b[58525] == 58525 && 
b[58526] == 58526 && 
b[58527] == 58527 && 
b[58528] == 58528 && 
b[58529] == 58529 && 
b[58530] == 58530 && 
b[58531] == 58531 && 
b[58532] == 58532 && 
b[58533] == 58533 && 
b[58534] == 58534 && 
b[58535] == 58535 && 
b[58536] == 58536 && 
b[58537] == 58537 && 
b[58538] == 58538 && 
b[58539] == 58539 && 
b[58540] == 58540 && 
b[58541] == 58541 && 
b[58542] == 58542 && 
b[58543] == 58543 && 
b[58544] == 58544 && 
b[58545] == 58545 && 
b[58546] == 58546 && 
b[58547] == 58547 && 
b[58548] == 58548 && 
b[58549] == 58549 && 
b[58550] == 58550 && 
b[58551] == 58551 && 
b[58552] == 58552 && 
b[58553] == 58553 && 
b[58554] == 58554 && 
b[58555] == 58555 && 
b[58556] == 58556 && 
b[58557] == 58557 && 
b[58558] == 58558 && 
b[58559] == 58559 && 
b[58560] == 58560 && 
b[58561] == 58561 && 
b[58562] == 58562 && 
b[58563] == 58563 && 
b[58564] == 58564 && 
b[58565] == 58565 && 
b[58566] == 58566 && 
b[58567] == 58567 && 
b[58568] == 58568 && 
b[58569] == 58569 && 
b[58570] == 58570 && 
b[58571] == 58571 && 
b[58572] == 58572 && 
b[58573] == 58573 && 
b[58574] == 58574 && 
b[58575] == 58575 && 
b[58576] == 58576 && 
b[58577] == 58577 && 
b[58578] == 58578 && 
b[58579] == 58579 && 
b[58580] == 58580 && 
b[58581] == 58581 && 
b[58582] == 58582 && 
b[58583] == 58583 && 
b[58584] == 58584 && 
b[58585] == 58585 && 
b[58586] == 58586 && 
b[58587] == 58587 && 
b[58588] == 58588 && 
b[58589] == 58589 && 
b[58590] == 58590 && 
b[58591] == 58591 && 
b[58592] == 58592 && 
b[58593] == 58593 && 
b[58594] == 58594 && 
b[58595] == 58595 && 
b[58596] == 58596 && 
b[58597] == 58597 && 
b[58598] == 58598 && 
b[58599] == 58599 && 
b[58600] == 58600 && 
b[58601] == 58601 && 
b[58602] == 58602 && 
b[58603] == 58603 && 
b[58604] == 58604 && 
b[58605] == 58605 && 
b[58606] == 58606 && 
b[58607] == 58607 && 
b[58608] == 58608 && 
b[58609] == 58609 && 
b[58610] == 58610 && 
b[58611] == 58611 && 
b[58612] == 58612 && 
b[58613] == 58613 && 
b[58614] == 58614 && 
b[58615] == 58615 && 
b[58616] == 58616 && 
b[58617] == 58617 && 
b[58618] == 58618 && 
b[58619] == 58619 && 
b[58620] == 58620 && 
b[58621] == 58621 && 
b[58622] == 58622 && 
b[58623] == 58623 && 
b[58624] == 58624 && 
b[58625] == 58625 && 
b[58626] == 58626 && 
b[58627] == 58627 && 
b[58628] == 58628 && 
b[58629] == 58629 && 
b[58630] == 58630 && 
b[58631] == 58631 && 
b[58632] == 58632 && 
b[58633] == 58633 && 
b[58634] == 58634 && 
b[58635] == 58635 && 
b[58636] == 58636 && 
b[58637] == 58637 && 
b[58638] == 58638 && 
b[58639] == 58639 && 
b[58640] == 58640 && 
b[58641] == 58641 && 
b[58642] == 58642 && 
b[58643] == 58643 && 
b[58644] == 58644 && 
b[58645] == 58645 && 
b[58646] == 58646 && 
b[58647] == 58647 && 
b[58648] == 58648 && 
b[58649] == 58649 && 
b[58650] == 58650 && 
b[58651] == 58651 && 
b[58652] == 58652 && 
b[58653] == 58653 && 
b[58654] == 58654 && 
b[58655] == 58655 && 
b[58656] == 58656 && 
b[58657] == 58657 && 
b[58658] == 58658 && 
b[58659] == 58659 && 
b[58660] == 58660 && 
b[58661] == 58661 && 
b[58662] == 58662 && 
b[58663] == 58663 && 
b[58664] == 58664 && 
b[58665] == 58665 && 
b[58666] == 58666 && 
b[58667] == 58667 && 
b[58668] == 58668 && 
b[58669] == 58669 && 
b[58670] == 58670 && 
b[58671] == 58671 && 
b[58672] == 58672 && 
b[58673] == 58673 && 
b[58674] == 58674 && 
b[58675] == 58675 && 
b[58676] == 58676 && 
b[58677] == 58677 && 
b[58678] == 58678 && 
b[58679] == 58679 && 
b[58680] == 58680 && 
b[58681] == 58681 && 
b[58682] == 58682 && 
b[58683] == 58683 && 
b[58684] == 58684 && 
b[58685] == 58685 && 
b[58686] == 58686 && 
b[58687] == 58687 && 
b[58688] == 58688 && 
b[58689] == 58689 && 
b[58690] == 58690 && 
b[58691] == 58691 && 
b[58692] == 58692 && 
b[58693] == 58693 && 
b[58694] == 58694 && 
b[58695] == 58695 && 
b[58696] == 58696 && 
b[58697] == 58697 && 
b[58698] == 58698 && 
b[58699] == 58699 && 
b[58700] == 58700 && 
b[58701] == 58701 && 
b[58702] == 58702 && 
b[58703] == 58703 && 
b[58704] == 58704 && 
b[58705] == 58705 && 
b[58706] == 58706 && 
b[58707] == 58707 && 
b[58708] == 58708 && 
b[58709] == 58709 && 
b[58710] == 58710 && 
b[58711] == 58711 && 
b[58712] == 58712 && 
b[58713] == 58713 && 
b[58714] == 58714 && 
b[58715] == 58715 && 
b[58716] == 58716 && 
b[58717] == 58717 && 
b[58718] == 58718 && 
b[58719] == 58719 && 
b[58720] == 58720 && 
b[58721] == 58721 && 
b[58722] == 58722 && 
b[58723] == 58723 && 
b[58724] == 58724 && 
b[58725] == 58725 && 
b[58726] == 58726 && 
b[58727] == 58727 && 
b[58728] == 58728 && 
b[58729] == 58729 && 
b[58730] == 58730 && 
b[58731] == 58731 && 
b[58732] == 58732 && 
b[58733] == 58733 && 
b[58734] == 58734 && 
b[58735] == 58735 && 
b[58736] == 58736 && 
b[58737] == 58737 && 
b[58738] == 58738 && 
b[58739] == 58739 && 
b[58740] == 58740 && 
b[58741] == 58741 && 
b[58742] == 58742 && 
b[58743] == 58743 && 
b[58744] == 58744 && 
b[58745] == 58745 && 
b[58746] == 58746 && 
b[58747] == 58747 && 
b[58748] == 58748 && 
b[58749] == 58749 && 
b[58750] == 58750 && 
b[58751] == 58751 && 
b[58752] == 58752 && 
b[58753] == 58753 && 
b[58754] == 58754 && 
b[58755] == 58755 && 
b[58756] == 58756 && 
b[58757] == 58757 && 
b[58758] == 58758 && 
b[58759] == 58759 && 
b[58760] == 58760 && 
b[58761] == 58761 && 
b[58762] == 58762 && 
b[58763] == 58763 && 
b[58764] == 58764 && 
b[58765] == 58765 && 
b[58766] == 58766 && 
b[58767] == 58767 && 
b[58768] == 58768 && 
b[58769] == 58769 && 
b[58770] == 58770 && 
b[58771] == 58771 && 
b[58772] == 58772 && 
b[58773] == 58773 && 
b[58774] == 58774 && 
b[58775] == 58775 && 
b[58776] == 58776 && 
b[58777] == 58777 && 
b[58778] == 58778 && 
b[58779] == 58779 && 
b[58780] == 58780 && 
b[58781] == 58781 && 
b[58782] == 58782 && 
b[58783] == 58783 && 
b[58784] == 58784 && 
b[58785] == 58785 && 
b[58786] == 58786 && 
b[58787] == 58787 && 
b[58788] == 58788 && 
b[58789] == 58789 && 
b[58790] == 58790 && 
b[58791] == 58791 && 
b[58792] == 58792 && 
b[58793] == 58793 && 
b[58794] == 58794 && 
b[58795] == 58795 && 
b[58796] == 58796 && 
b[58797] == 58797 && 
b[58798] == 58798 && 
b[58799] == 58799 && 
b[58800] == 58800 && 
b[58801] == 58801 && 
b[58802] == 58802 && 
b[58803] == 58803 && 
b[58804] == 58804 && 
b[58805] == 58805 && 
b[58806] == 58806 && 
b[58807] == 58807 && 
b[58808] == 58808 && 
b[58809] == 58809 && 
b[58810] == 58810 && 
b[58811] == 58811 && 
b[58812] == 58812 && 
b[58813] == 58813 && 
b[58814] == 58814 && 
b[58815] == 58815 && 
b[58816] == 58816 && 
b[58817] == 58817 && 
b[58818] == 58818 && 
b[58819] == 58819 && 
b[58820] == 58820 && 
b[58821] == 58821 && 
b[58822] == 58822 && 
b[58823] == 58823 && 
b[58824] == 58824 && 
b[58825] == 58825 && 
b[58826] == 58826 && 
b[58827] == 58827 && 
b[58828] == 58828 && 
b[58829] == 58829 && 
b[58830] == 58830 && 
b[58831] == 58831 && 
b[58832] == 58832 && 
b[58833] == 58833 && 
b[58834] == 58834 && 
b[58835] == 58835 && 
b[58836] == 58836 && 
b[58837] == 58837 && 
b[58838] == 58838 && 
b[58839] == 58839 && 
b[58840] == 58840 && 
b[58841] == 58841 && 
b[58842] == 58842 && 
b[58843] == 58843 && 
b[58844] == 58844 && 
b[58845] == 58845 && 
b[58846] == 58846 && 
b[58847] == 58847 && 
b[58848] == 58848 && 
b[58849] == 58849 && 
b[58850] == 58850 && 
b[58851] == 58851 && 
b[58852] == 58852 && 
b[58853] == 58853 && 
b[58854] == 58854 && 
b[58855] == 58855 && 
b[58856] == 58856 && 
b[58857] == 58857 && 
b[58858] == 58858 && 
b[58859] == 58859 && 
b[58860] == 58860 && 
b[58861] == 58861 && 
b[58862] == 58862 && 
b[58863] == 58863 && 
b[58864] == 58864 && 
b[58865] == 58865 && 
b[58866] == 58866 && 
b[58867] == 58867 && 
b[58868] == 58868 && 
b[58869] == 58869 && 
b[58870] == 58870 && 
b[58871] == 58871 && 
b[58872] == 58872 && 
b[58873] == 58873 && 
b[58874] == 58874 && 
b[58875] == 58875 && 
b[58876] == 58876 && 
b[58877] == 58877 && 
b[58878] == 58878 && 
b[58879] == 58879 && 
b[58880] == 58880 && 
b[58881] == 58881 && 
b[58882] == 58882 && 
b[58883] == 58883 && 
b[58884] == 58884 && 
b[58885] == 58885 && 
b[58886] == 58886 && 
b[58887] == 58887 && 
b[58888] == 58888 && 
b[58889] == 58889 && 
b[58890] == 58890 && 
b[58891] == 58891 && 
b[58892] == 58892 && 
b[58893] == 58893 && 
b[58894] == 58894 && 
b[58895] == 58895 && 
b[58896] == 58896 && 
b[58897] == 58897 && 
b[58898] == 58898 && 
b[58899] == 58899 && 
b[58900] == 58900 && 
b[58901] == 58901 && 
b[58902] == 58902 && 
b[58903] == 58903 && 
b[58904] == 58904 && 
b[58905] == 58905 && 
b[58906] == 58906 && 
b[58907] == 58907 && 
b[58908] == 58908 && 
b[58909] == 58909 && 
b[58910] == 58910 && 
b[58911] == 58911 && 
b[58912] == 58912 && 
b[58913] == 58913 && 
b[58914] == 58914 && 
b[58915] == 58915 && 
b[58916] == 58916 && 
b[58917] == 58917 && 
b[58918] == 58918 && 
b[58919] == 58919 && 
b[58920] == 58920 && 
b[58921] == 58921 && 
b[58922] == 58922 && 
b[58923] == 58923 && 
b[58924] == 58924 && 
b[58925] == 58925 && 
b[58926] == 58926 && 
b[58927] == 58927 && 
b[58928] == 58928 && 
b[58929] == 58929 && 
b[58930] == 58930 && 
b[58931] == 58931 && 
b[58932] == 58932 && 
b[58933] == 58933 && 
b[58934] == 58934 && 
b[58935] == 58935 && 
b[58936] == 58936 && 
b[58937] == 58937 && 
b[58938] == 58938 && 
b[58939] == 58939 && 
b[58940] == 58940 && 
b[58941] == 58941 && 
b[58942] == 58942 && 
b[58943] == 58943 && 
b[58944] == 58944 && 
b[58945] == 58945 && 
b[58946] == 58946 && 
b[58947] == 58947 && 
b[58948] == 58948 && 
b[58949] == 58949 && 
b[58950] == 58950 && 
b[58951] == 58951 && 
b[58952] == 58952 && 
b[58953] == 58953 && 
b[58954] == 58954 && 
b[58955] == 58955 && 
b[58956] == 58956 && 
b[58957] == 58957 && 
b[58958] == 58958 && 
b[58959] == 58959 && 
b[58960] == 58960 && 
b[58961] == 58961 && 
b[58962] == 58962 && 
b[58963] == 58963 && 
b[58964] == 58964 && 
b[58965] == 58965 && 
b[58966] == 58966 && 
b[58967] == 58967 && 
b[58968] == 58968 && 
b[58969] == 58969 && 
b[58970] == 58970 && 
b[58971] == 58971 && 
b[58972] == 58972 && 
b[58973] == 58973 && 
b[58974] == 58974 && 
b[58975] == 58975 && 
b[58976] == 58976 && 
b[58977] == 58977 && 
b[58978] == 58978 && 
b[58979] == 58979 && 
b[58980] == 58980 && 
b[58981] == 58981 && 
b[58982] == 58982 && 
b[58983] == 58983 && 
b[58984] == 58984 && 
b[58985] == 58985 && 
b[58986] == 58986 && 
b[58987] == 58987 && 
b[58988] == 58988 && 
b[58989] == 58989 && 
b[58990] == 58990 && 
b[58991] == 58991 && 
b[58992] == 58992 && 
b[58993] == 58993 && 
b[58994] == 58994 && 
b[58995] == 58995 && 
b[58996] == 58996 && 
b[58997] == 58997 && 
b[58998] == 58998 && 
b[58999] == 58999 && 
b[59000] == 59000 && 
b[59001] == 59001 && 
b[59002] == 59002 && 
b[59003] == 59003 && 
b[59004] == 59004 && 
b[59005] == 59005 && 
b[59006] == 59006 && 
b[59007] == 59007 && 
b[59008] == 59008 && 
b[59009] == 59009 && 
b[59010] == 59010 && 
b[59011] == 59011 && 
b[59012] == 59012 && 
b[59013] == 59013 && 
b[59014] == 59014 && 
b[59015] == 59015 && 
b[59016] == 59016 && 
b[59017] == 59017 && 
b[59018] == 59018 && 
b[59019] == 59019 && 
b[59020] == 59020 && 
b[59021] == 59021 && 
b[59022] == 59022 && 
b[59023] == 59023 && 
b[59024] == 59024 && 
b[59025] == 59025 && 
b[59026] == 59026 && 
b[59027] == 59027 && 
b[59028] == 59028 && 
b[59029] == 59029 && 
b[59030] == 59030 && 
b[59031] == 59031 && 
b[59032] == 59032 && 
b[59033] == 59033 && 
b[59034] == 59034 && 
b[59035] == 59035 && 
b[59036] == 59036 && 
b[59037] == 59037 && 
b[59038] == 59038 && 
b[59039] == 59039 && 
b[59040] == 59040 && 
b[59041] == 59041 && 
b[59042] == 59042 && 
b[59043] == 59043 && 
b[59044] == 59044 && 
b[59045] == 59045 && 
b[59046] == 59046 && 
b[59047] == 59047 && 
b[59048] == 59048 && 
b[59049] == 59049 && 
b[59050] == 59050 && 
b[59051] == 59051 && 
b[59052] == 59052 && 
b[59053] == 59053 && 
b[59054] == 59054 && 
b[59055] == 59055 && 
b[59056] == 59056 && 
b[59057] == 59057 && 
b[59058] == 59058 && 
b[59059] == 59059 && 
b[59060] == 59060 && 
b[59061] == 59061 && 
b[59062] == 59062 && 
b[59063] == 59063 && 
b[59064] == 59064 && 
b[59065] == 59065 && 
b[59066] == 59066 && 
b[59067] == 59067 && 
b[59068] == 59068 && 
b[59069] == 59069 && 
b[59070] == 59070 && 
b[59071] == 59071 && 
b[59072] == 59072 && 
b[59073] == 59073 && 
b[59074] == 59074 && 
b[59075] == 59075 && 
b[59076] == 59076 && 
b[59077] == 59077 && 
b[59078] == 59078 && 
b[59079] == 59079 && 
b[59080] == 59080 && 
b[59081] == 59081 && 
b[59082] == 59082 && 
b[59083] == 59083 && 
b[59084] == 59084 && 
b[59085] == 59085 && 
b[59086] == 59086 && 
b[59087] == 59087 && 
b[59088] == 59088 && 
b[59089] == 59089 && 
b[59090] == 59090 && 
b[59091] == 59091 && 
b[59092] == 59092 && 
b[59093] == 59093 && 
b[59094] == 59094 && 
b[59095] == 59095 && 
b[59096] == 59096 && 
b[59097] == 59097 && 
b[59098] == 59098 && 
b[59099] == 59099 && 
b[59100] == 59100 && 
b[59101] == 59101 && 
b[59102] == 59102 && 
b[59103] == 59103 && 
b[59104] == 59104 && 
b[59105] == 59105 && 
b[59106] == 59106 && 
b[59107] == 59107 && 
b[59108] == 59108 && 
b[59109] == 59109 && 
b[59110] == 59110 && 
b[59111] == 59111 && 
b[59112] == 59112 && 
b[59113] == 59113 && 
b[59114] == 59114 && 
b[59115] == 59115 && 
b[59116] == 59116 && 
b[59117] == 59117 && 
b[59118] == 59118 && 
b[59119] == 59119 && 
b[59120] == 59120 && 
b[59121] == 59121 && 
b[59122] == 59122 && 
b[59123] == 59123 && 
b[59124] == 59124 && 
b[59125] == 59125 && 
b[59126] == 59126 && 
b[59127] == 59127 && 
b[59128] == 59128 && 
b[59129] == 59129 && 
b[59130] == 59130 && 
b[59131] == 59131 && 
b[59132] == 59132 && 
b[59133] == 59133 && 
b[59134] == 59134 && 
b[59135] == 59135 && 
b[59136] == 59136 && 
b[59137] == 59137 && 
b[59138] == 59138 && 
b[59139] == 59139 && 
b[59140] == 59140 && 
b[59141] == 59141 && 
b[59142] == 59142 && 
b[59143] == 59143 && 
b[59144] == 59144 && 
b[59145] == 59145 && 
b[59146] == 59146 && 
b[59147] == 59147 && 
b[59148] == 59148 && 
b[59149] == 59149 && 
b[59150] == 59150 && 
b[59151] == 59151 && 
b[59152] == 59152 && 
b[59153] == 59153 && 
b[59154] == 59154 && 
b[59155] == 59155 && 
b[59156] == 59156 && 
b[59157] == 59157 && 
b[59158] == 59158 && 
b[59159] == 59159 && 
b[59160] == 59160 && 
b[59161] == 59161 && 
b[59162] == 59162 && 
b[59163] == 59163 && 
b[59164] == 59164 && 
b[59165] == 59165 && 
b[59166] == 59166 && 
b[59167] == 59167 && 
b[59168] == 59168 && 
b[59169] == 59169 && 
b[59170] == 59170 && 
b[59171] == 59171 && 
b[59172] == 59172 && 
b[59173] == 59173 && 
b[59174] == 59174 && 
b[59175] == 59175 && 
b[59176] == 59176 && 
b[59177] == 59177 && 
b[59178] == 59178 && 
b[59179] == 59179 && 
b[59180] == 59180 && 
b[59181] == 59181 && 
b[59182] == 59182 && 
b[59183] == 59183 && 
b[59184] == 59184 && 
b[59185] == 59185 && 
b[59186] == 59186 && 
b[59187] == 59187 && 
b[59188] == 59188 && 
b[59189] == 59189 && 
b[59190] == 59190 && 
b[59191] == 59191 && 
b[59192] == 59192 && 
b[59193] == 59193 && 
b[59194] == 59194 && 
b[59195] == 59195 && 
b[59196] == 59196 && 
b[59197] == 59197 && 
b[59198] == 59198 && 
b[59199] == 59199 && 
b[59200] == 59200 && 
b[59201] == 59201 && 
b[59202] == 59202 && 
b[59203] == 59203 && 
b[59204] == 59204 && 
b[59205] == 59205 && 
b[59206] == 59206 && 
b[59207] == 59207 && 
b[59208] == 59208 && 
b[59209] == 59209 && 
b[59210] == 59210 && 
b[59211] == 59211 && 
b[59212] == 59212 && 
b[59213] == 59213 && 
b[59214] == 59214 && 
b[59215] == 59215 && 
b[59216] == 59216 && 
b[59217] == 59217 && 
b[59218] == 59218 && 
b[59219] == 59219 && 
b[59220] == 59220 && 
b[59221] == 59221 && 
b[59222] == 59222 && 
b[59223] == 59223 && 
b[59224] == 59224 && 
b[59225] == 59225 && 
b[59226] == 59226 && 
b[59227] == 59227 && 
b[59228] == 59228 && 
b[59229] == 59229 && 
b[59230] == 59230 && 
b[59231] == 59231 && 
b[59232] == 59232 && 
b[59233] == 59233 && 
b[59234] == 59234 && 
b[59235] == 59235 && 
b[59236] == 59236 && 
b[59237] == 59237 && 
b[59238] == 59238 && 
b[59239] == 59239 && 
b[59240] == 59240 && 
b[59241] == 59241 && 
b[59242] == 59242 && 
b[59243] == 59243 && 
b[59244] == 59244 && 
b[59245] == 59245 && 
b[59246] == 59246 && 
b[59247] == 59247 && 
b[59248] == 59248 && 
b[59249] == 59249 && 
b[59250] == 59250 && 
b[59251] == 59251 && 
b[59252] == 59252 && 
b[59253] == 59253 && 
b[59254] == 59254 && 
b[59255] == 59255 && 
b[59256] == 59256 && 
b[59257] == 59257 && 
b[59258] == 59258 && 
b[59259] == 59259 && 
b[59260] == 59260 && 
b[59261] == 59261 && 
b[59262] == 59262 && 
b[59263] == 59263 && 
b[59264] == 59264 && 
b[59265] == 59265 && 
b[59266] == 59266 && 
b[59267] == 59267 && 
b[59268] == 59268 && 
b[59269] == 59269 && 
b[59270] == 59270 && 
b[59271] == 59271 && 
b[59272] == 59272 && 
b[59273] == 59273 && 
b[59274] == 59274 && 
b[59275] == 59275 && 
b[59276] == 59276 && 
b[59277] == 59277 && 
b[59278] == 59278 && 
b[59279] == 59279 && 
b[59280] == 59280 && 
b[59281] == 59281 && 
b[59282] == 59282 && 
b[59283] == 59283 && 
b[59284] == 59284 && 
b[59285] == 59285 && 
b[59286] == 59286 && 
b[59287] == 59287 && 
b[59288] == 59288 && 
b[59289] == 59289 && 
b[59290] == 59290 && 
b[59291] == 59291 && 
b[59292] == 59292 && 
b[59293] == 59293 && 
b[59294] == 59294 && 
b[59295] == 59295 && 
b[59296] == 59296 && 
b[59297] == 59297 && 
b[59298] == 59298 && 
b[59299] == 59299 && 
b[59300] == 59300 && 
b[59301] == 59301 && 
b[59302] == 59302 && 
b[59303] == 59303 && 
b[59304] == 59304 && 
b[59305] == 59305 && 
b[59306] == 59306 && 
b[59307] == 59307 && 
b[59308] == 59308 && 
b[59309] == 59309 && 
b[59310] == 59310 && 
b[59311] == 59311 && 
b[59312] == 59312 && 
b[59313] == 59313 && 
b[59314] == 59314 && 
b[59315] == 59315 && 
b[59316] == 59316 && 
b[59317] == 59317 && 
b[59318] == 59318 && 
b[59319] == 59319 && 
b[59320] == 59320 && 
b[59321] == 59321 && 
b[59322] == 59322 && 
b[59323] == 59323 && 
b[59324] == 59324 && 
b[59325] == 59325 && 
b[59326] == 59326 && 
b[59327] == 59327 && 
b[59328] == 59328 && 
b[59329] == 59329 && 
b[59330] == 59330 && 
b[59331] == 59331 && 
b[59332] == 59332 && 
b[59333] == 59333 && 
b[59334] == 59334 && 
b[59335] == 59335 && 
b[59336] == 59336 && 
b[59337] == 59337 && 
b[59338] == 59338 && 
b[59339] == 59339 && 
b[59340] == 59340 && 
b[59341] == 59341 && 
b[59342] == 59342 && 
b[59343] == 59343 && 
b[59344] == 59344 && 
b[59345] == 59345 && 
b[59346] == 59346 && 
b[59347] == 59347 && 
b[59348] == 59348 && 
b[59349] == 59349 && 
b[59350] == 59350 && 
b[59351] == 59351 && 
b[59352] == 59352 && 
b[59353] == 59353 && 
b[59354] == 59354 && 
b[59355] == 59355 && 
b[59356] == 59356 && 
b[59357] == 59357 && 
b[59358] == 59358 && 
b[59359] == 59359 && 
b[59360] == 59360 && 
b[59361] == 59361 && 
b[59362] == 59362 && 
b[59363] == 59363 && 
b[59364] == 59364 && 
b[59365] == 59365 && 
b[59366] == 59366 && 
b[59367] == 59367 && 
b[59368] == 59368 && 
b[59369] == 59369 && 
b[59370] == 59370 && 
b[59371] == 59371 && 
b[59372] == 59372 && 
b[59373] == 59373 && 
b[59374] == 59374 && 
b[59375] == 59375 && 
b[59376] == 59376 && 
b[59377] == 59377 && 
b[59378] == 59378 && 
b[59379] == 59379 && 
b[59380] == 59380 && 
b[59381] == 59381 && 
b[59382] == 59382 && 
b[59383] == 59383 && 
b[59384] == 59384 && 
b[59385] == 59385 && 
b[59386] == 59386 && 
b[59387] == 59387 && 
b[59388] == 59388 && 
b[59389] == 59389 && 
b[59390] == 59390 && 
b[59391] == 59391 && 
b[59392] == 59392 && 
b[59393] == 59393 && 
b[59394] == 59394 && 
b[59395] == 59395 && 
b[59396] == 59396 && 
b[59397] == 59397 && 
b[59398] == 59398 && 
b[59399] == 59399 && 
b[59400] == 59400 && 
b[59401] == 59401 && 
b[59402] == 59402 && 
b[59403] == 59403 && 
b[59404] == 59404 && 
b[59405] == 59405 && 
b[59406] == 59406 && 
b[59407] == 59407 && 
b[59408] == 59408 && 
b[59409] == 59409 && 
b[59410] == 59410 && 
b[59411] == 59411 && 
b[59412] == 59412 && 
b[59413] == 59413 && 
b[59414] == 59414 && 
b[59415] == 59415 && 
b[59416] == 59416 && 
b[59417] == 59417 && 
b[59418] == 59418 && 
b[59419] == 59419 && 
b[59420] == 59420 && 
b[59421] == 59421 && 
b[59422] == 59422 && 
b[59423] == 59423 && 
b[59424] == 59424 && 
b[59425] == 59425 && 
b[59426] == 59426 && 
b[59427] == 59427 && 
b[59428] == 59428 && 
b[59429] == 59429 && 
b[59430] == 59430 && 
b[59431] == 59431 && 
b[59432] == 59432 && 
b[59433] == 59433 && 
b[59434] == 59434 && 
b[59435] == 59435 && 
b[59436] == 59436 && 
b[59437] == 59437 && 
b[59438] == 59438 && 
b[59439] == 59439 && 
b[59440] == 59440 && 
b[59441] == 59441 && 
b[59442] == 59442 && 
b[59443] == 59443 && 
b[59444] == 59444 && 
b[59445] == 59445 && 
b[59446] == 59446 && 
b[59447] == 59447 && 
b[59448] == 59448 && 
b[59449] == 59449 && 
b[59450] == 59450 && 
b[59451] == 59451 && 
b[59452] == 59452 && 
b[59453] == 59453 && 
b[59454] == 59454 && 
b[59455] == 59455 && 
b[59456] == 59456 && 
b[59457] == 59457 && 
b[59458] == 59458 && 
b[59459] == 59459 && 
b[59460] == 59460 && 
b[59461] == 59461 && 
b[59462] == 59462 && 
b[59463] == 59463 && 
b[59464] == 59464 && 
b[59465] == 59465 && 
b[59466] == 59466 && 
b[59467] == 59467 && 
b[59468] == 59468 && 
b[59469] == 59469 && 
b[59470] == 59470 && 
b[59471] == 59471 && 
b[59472] == 59472 && 
b[59473] == 59473 && 
b[59474] == 59474 && 
b[59475] == 59475 && 
b[59476] == 59476 && 
b[59477] == 59477 && 
b[59478] == 59478 && 
b[59479] == 59479 && 
b[59480] == 59480 && 
b[59481] == 59481 && 
b[59482] == 59482 && 
b[59483] == 59483 && 
b[59484] == 59484 && 
b[59485] == 59485 && 
b[59486] == 59486 && 
b[59487] == 59487 && 
b[59488] == 59488 && 
b[59489] == 59489 && 
b[59490] == 59490 && 
b[59491] == 59491 && 
b[59492] == 59492 && 
b[59493] == 59493 && 
b[59494] == 59494 && 
b[59495] == 59495 && 
b[59496] == 59496 && 
b[59497] == 59497 && 
b[59498] == 59498 && 
b[59499] == 59499 && 
b[59500] == 59500 && 
b[59501] == 59501 && 
b[59502] == 59502 && 
b[59503] == 59503 && 
b[59504] == 59504 && 
b[59505] == 59505 && 
b[59506] == 59506 && 
b[59507] == 59507 && 
b[59508] == 59508 && 
b[59509] == 59509 && 
b[59510] == 59510 && 
b[59511] == 59511 && 
b[59512] == 59512 && 
b[59513] == 59513 && 
b[59514] == 59514 && 
b[59515] == 59515 && 
b[59516] == 59516 && 
b[59517] == 59517 && 
b[59518] == 59518 && 
b[59519] == 59519 && 
b[59520] == 59520 && 
b[59521] == 59521 && 
b[59522] == 59522 && 
b[59523] == 59523 && 
b[59524] == 59524 && 
b[59525] == 59525 && 
b[59526] == 59526 && 
b[59527] == 59527 && 
b[59528] == 59528 && 
b[59529] == 59529 && 
b[59530] == 59530 && 
b[59531] == 59531 && 
b[59532] == 59532 && 
b[59533] == 59533 && 
b[59534] == 59534 && 
b[59535] == 59535 && 
b[59536] == 59536 && 
b[59537] == 59537 && 
b[59538] == 59538 && 
b[59539] == 59539 && 
b[59540] == 59540 && 
b[59541] == 59541 && 
b[59542] == 59542 && 
b[59543] == 59543 && 
b[59544] == 59544 && 
b[59545] == 59545 && 
b[59546] == 59546 && 
b[59547] == 59547 && 
b[59548] == 59548 && 
b[59549] == 59549 && 
b[59550] == 59550 && 
b[59551] == 59551 && 
b[59552] == 59552 && 
b[59553] == 59553 && 
b[59554] == 59554 && 
b[59555] == 59555 && 
b[59556] == 59556 && 
b[59557] == 59557 && 
b[59558] == 59558 && 
b[59559] == 59559 && 
b[59560] == 59560 && 
b[59561] == 59561 && 
b[59562] == 59562 && 
b[59563] == 59563 && 
b[59564] == 59564 && 
b[59565] == 59565 && 
b[59566] == 59566 && 
b[59567] == 59567 && 
b[59568] == 59568 && 
b[59569] == 59569 && 
b[59570] == 59570 && 
b[59571] == 59571 && 
b[59572] == 59572 && 
b[59573] == 59573 && 
b[59574] == 59574 && 
b[59575] == 59575 && 
b[59576] == 59576 && 
b[59577] == 59577 && 
b[59578] == 59578 && 
b[59579] == 59579 && 
b[59580] == 59580 && 
b[59581] == 59581 && 
b[59582] == 59582 && 
b[59583] == 59583 && 
b[59584] == 59584 && 
b[59585] == 59585 && 
b[59586] == 59586 && 
b[59587] == 59587 && 
b[59588] == 59588 && 
b[59589] == 59589 && 
b[59590] == 59590 && 
b[59591] == 59591 && 
b[59592] == 59592 && 
b[59593] == 59593 && 
b[59594] == 59594 && 
b[59595] == 59595 && 
b[59596] == 59596 && 
b[59597] == 59597 && 
b[59598] == 59598 && 
b[59599] == 59599 && 
b[59600] == 59600 && 
b[59601] == 59601 && 
b[59602] == 59602 && 
b[59603] == 59603 && 
b[59604] == 59604 && 
b[59605] == 59605 && 
b[59606] == 59606 && 
b[59607] == 59607 && 
b[59608] == 59608 && 
b[59609] == 59609 && 
b[59610] == 59610 && 
b[59611] == 59611 && 
b[59612] == 59612 && 
b[59613] == 59613 && 
b[59614] == 59614 && 
b[59615] == 59615 && 
b[59616] == 59616 && 
b[59617] == 59617 && 
b[59618] == 59618 && 
b[59619] == 59619 && 
b[59620] == 59620 && 
b[59621] == 59621 && 
b[59622] == 59622 && 
b[59623] == 59623 && 
b[59624] == 59624 && 
b[59625] == 59625 && 
b[59626] == 59626 && 
b[59627] == 59627 && 
b[59628] == 59628 && 
b[59629] == 59629 && 
b[59630] == 59630 && 
b[59631] == 59631 && 
b[59632] == 59632 && 
b[59633] == 59633 && 
b[59634] == 59634 && 
b[59635] == 59635 && 
b[59636] == 59636 && 
b[59637] == 59637 && 
b[59638] == 59638 && 
b[59639] == 59639 && 
b[59640] == 59640 && 
b[59641] == 59641 && 
b[59642] == 59642 && 
b[59643] == 59643 && 
b[59644] == 59644 && 
b[59645] == 59645 && 
b[59646] == 59646 && 
b[59647] == 59647 && 
b[59648] == 59648 && 
b[59649] == 59649 && 
b[59650] == 59650 && 
b[59651] == 59651 && 
b[59652] == 59652 && 
b[59653] == 59653 && 
b[59654] == 59654 && 
b[59655] == 59655 && 
b[59656] == 59656 && 
b[59657] == 59657 && 
b[59658] == 59658 && 
b[59659] == 59659 && 
b[59660] == 59660 && 
b[59661] == 59661 && 
b[59662] == 59662 && 
b[59663] == 59663 && 
b[59664] == 59664 && 
b[59665] == 59665 && 
b[59666] == 59666 && 
b[59667] == 59667 && 
b[59668] == 59668 && 
b[59669] == 59669 && 
b[59670] == 59670 && 
b[59671] == 59671 && 
b[59672] == 59672 && 
b[59673] == 59673 && 
b[59674] == 59674 && 
b[59675] == 59675 && 
b[59676] == 59676 && 
b[59677] == 59677 && 
b[59678] == 59678 && 
b[59679] == 59679 && 
b[59680] == 59680 && 
b[59681] == 59681 && 
b[59682] == 59682 && 
b[59683] == 59683 && 
b[59684] == 59684 && 
b[59685] == 59685 && 
b[59686] == 59686 && 
b[59687] == 59687 && 
b[59688] == 59688 && 
b[59689] == 59689 && 
b[59690] == 59690 && 
b[59691] == 59691 && 
b[59692] == 59692 && 
b[59693] == 59693 && 
b[59694] == 59694 && 
b[59695] == 59695 && 
b[59696] == 59696 && 
b[59697] == 59697 && 
b[59698] == 59698 && 
b[59699] == 59699 && 
b[59700] == 59700 && 
b[59701] == 59701 && 
b[59702] == 59702 && 
b[59703] == 59703 && 
b[59704] == 59704 && 
b[59705] == 59705 && 
b[59706] == 59706 && 
b[59707] == 59707 && 
b[59708] == 59708 && 
b[59709] == 59709 && 
b[59710] == 59710 && 
b[59711] == 59711 && 
b[59712] == 59712 && 
b[59713] == 59713 && 
b[59714] == 59714 && 
b[59715] == 59715 && 
b[59716] == 59716 && 
b[59717] == 59717 && 
b[59718] == 59718 && 
b[59719] == 59719 && 
b[59720] == 59720 && 
b[59721] == 59721 && 
b[59722] == 59722 && 
b[59723] == 59723 && 
b[59724] == 59724 && 
b[59725] == 59725 && 
b[59726] == 59726 && 
b[59727] == 59727 && 
b[59728] == 59728 && 
b[59729] == 59729 && 
b[59730] == 59730 && 
b[59731] == 59731 && 
b[59732] == 59732 && 
b[59733] == 59733 && 
b[59734] == 59734 && 
b[59735] == 59735 && 
b[59736] == 59736 && 
b[59737] == 59737 && 
b[59738] == 59738 && 
b[59739] == 59739 && 
b[59740] == 59740 && 
b[59741] == 59741 && 
b[59742] == 59742 && 
b[59743] == 59743 && 
b[59744] == 59744 && 
b[59745] == 59745 && 
b[59746] == 59746 && 
b[59747] == 59747 && 
b[59748] == 59748 && 
b[59749] == 59749 && 
b[59750] == 59750 && 
b[59751] == 59751 && 
b[59752] == 59752 && 
b[59753] == 59753 && 
b[59754] == 59754 && 
b[59755] == 59755 && 
b[59756] == 59756 && 
b[59757] == 59757 && 
b[59758] == 59758 && 
b[59759] == 59759 && 
b[59760] == 59760 && 
b[59761] == 59761 && 
b[59762] == 59762 && 
b[59763] == 59763 && 
b[59764] == 59764 && 
b[59765] == 59765 && 
b[59766] == 59766 && 
b[59767] == 59767 && 
b[59768] == 59768 && 
b[59769] == 59769 && 
b[59770] == 59770 && 
b[59771] == 59771 && 
b[59772] == 59772 && 
b[59773] == 59773 && 
b[59774] == 59774 && 
b[59775] == 59775 && 
b[59776] == 59776 && 
b[59777] == 59777 && 
b[59778] == 59778 && 
b[59779] == 59779 && 
b[59780] == 59780 && 
b[59781] == 59781 && 
b[59782] == 59782 && 
b[59783] == 59783 && 
b[59784] == 59784 && 
b[59785] == 59785 && 
b[59786] == 59786 && 
b[59787] == 59787 && 
b[59788] == 59788 && 
b[59789] == 59789 && 
b[59790] == 59790 && 
b[59791] == 59791 && 
b[59792] == 59792 && 
b[59793] == 59793 && 
b[59794] == 59794 && 
b[59795] == 59795 && 
b[59796] == 59796 && 
b[59797] == 59797 && 
b[59798] == 59798 && 
b[59799] == 59799 && 
b[59800] == 59800 && 
b[59801] == 59801 && 
b[59802] == 59802 && 
b[59803] == 59803 && 
b[59804] == 59804 && 
b[59805] == 59805 && 
b[59806] == 59806 && 
b[59807] == 59807 && 
b[59808] == 59808 && 
b[59809] == 59809 && 
b[59810] == 59810 && 
b[59811] == 59811 && 
b[59812] == 59812 && 
b[59813] == 59813 && 
b[59814] == 59814 && 
b[59815] == 59815 && 
b[59816] == 59816 && 
b[59817] == 59817 && 
b[59818] == 59818 && 
b[59819] == 59819 && 
b[59820] == 59820 && 
b[59821] == 59821 && 
b[59822] == 59822 && 
b[59823] == 59823 && 
b[59824] == 59824 && 
b[59825] == 59825 && 
b[59826] == 59826 && 
b[59827] == 59827 && 
b[59828] == 59828 && 
b[59829] == 59829 && 
b[59830] == 59830 && 
b[59831] == 59831 && 
b[59832] == 59832 && 
b[59833] == 59833 && 
b[59834] == 59834 && 
b[59835] == 59835 && 
b[59836] == 59836 && 
b[59837] == 59837 && 
b[59838] == 59838 && 
b[59839] == 59839 && 
b[59840] == 59840 && 
b[59841] == 59841 && 
b[59842] == 59842 && 
b[59843] == 59843 && 
b[59844] == 59844 && 
b[59845] == 59845 && 
b[59846] == 59846 && 
b[59847] == 59847 && 
b[59848] == 59848 && 
b[59849] == 59849 && 
b[59850] == 59850 && 
b[59851] == 59851 && 
b[59852] == 59852 && 
b[59853] == 59853 && 
b[59854] == 59854 && 
b[59855] == 59855 && 
b[59856] == 59856 && 
b[59857] == 59857 && 
b[59858] == 59858 && 
b[59859] == 59859 && 
b[59860] == 59860 && 
b[59861] == 59861 && 
b[59862] == 59862 && 
b[59863] == 59863 && 
b[59864] == 59864 && 
b[59865] == 59865 && 
b[59866] == 59866 && 
b[59867] == 59867 && 
b[59868] == 59868 && 
b[59869] == 59869 && 
b[59870] == 59870 && 
b[59871] == 59871 && 
b[59872] == 59872 && 
b[59873] == 59873 && 
b[59874] == 59874 && 
b[59875] == 59875 && 
b[59876] == 59876 && 
b[59877] == 59877 && 
b[59878] == 59878 && 
b[59879] == 59879 && 
b[59880] == 59880 && 
b[59881] == 59881 && 
b[59882] == 59882 && 
b[59883] == 59883 && 
b[59884] == 59884 && 
b[59885] == 59885 && 
b[59886] == 59886 && 
b[59887] == 59887 && 
b[59888] == 59888 && 
b[59889] == 59889 && 
b[59890] == 59890 && 
b[59891] == 59891 && 
b[59892] == 59892 && 
b[59893] == 59893 && 
b[59894] == 59894 && 
b[59895] == 59895 && 
b[59896] == 59896 && 
b[59897] == 59897 && 
b[59898] == 59898 && 
b[59899] == 59899 && 
b[59900] == 59900 && 
b[59901] == 59901 && 
b[59902] == 59902 && 
b[59903] == 59903 && 
b[59904] == 59904 && 
b[59905] == 59905 && 
b[59906] == 59906 && 
b[59907] == 59907 && 
b[59908] == 59908 && 
b[59909] == 59909 && 
b[59910] == 59910 && 
b[59911] == 59911 && 
b[59912] == 59912 && 
b[59913] == 59913 && 
b[59914] == 59914 && 
b[59915] == 59915 && 
b[59916] == 59916 && 
b[59917] == 59917 && 
b[59918] == 59918 && 
b[59919] == 59919 && 
b[59920] == 59920 && 
b[59921] == 59921 && 
b[59922] == 59922 && 
b[59923] == 59923 && 
b[59924] == 59924 && 
b[59925] == 59925 && 
b[59926] == 59926 && 
b[59927] == 59927 && 
b[59928] == 59928 && 
b[59929] == 59929 && 
b[59930] == 59930 && 
b[59931] == 59931 && 
b[59932] == 59932 && 
b[59933] == 59933 && 
b[59934] == 59934 && 
b[59935] == 59935 && 
b[59936] == 59936 && 
b[59937] == 59937 && 
b[59938] == 59938 && 
b[59939] == 59939 && 
b[59940] == 59940 && 
b[59941] == 59941 && 
b[59942] == 59942 && 
b[59943] == 59943 && 
b[59944] == 59944 && 
b[59945] == 59945 && 
b[59946] == 59946 && 
b[59947] == 59947 && 
b[59948] == 59948 && 
b[59949] == 59949 && 
b[59950] == 59950 && 
b[59951] == 59951 && 
b[59952] == 59952 && 
b[59953] == 59953 && 
b[59954] == 59954 && 
b[59955] == 59955 && 
b[59956] == 59956 && 
b[59957] == 59957 && 
b[59958] == 59958 && 
b[59959] == 59959 && 
b[59960] == 59960 && 
b[59961] == 59961 && 
b[59962] == 59962 && 
b[59963] == 59963 && 
b[59964] == 59964 && 
b[59965] == 59965 && 
b[59966] == 59966 && 
b[59967] == 59967 && 
b[59968] == 59968 && 
b[59969] == 59969 && 
b[59970] == 59970 && 
b[59971] == 59971 && 
b[59972] == 59972 && 
b[59973] == 59973 && 
b[59974] == 59974 && 
b[59975] == 59975 && 
b[59976] == 59976 && 
b[59977] == 59977 && 
b[59978] == 59978 && 
b[59979] == 59979 && 
b[59980] == 59980 && 
b[59981] == 59981 && 
b[59982] == 59982 && 
b[59983] == 59983 && 
b[59984] == 59984 && 
b[59985] == 59985 && 
b[59986] == 59986 && 
b[59987] == 59987 && 
b[59988] == 59988 && 
b[59989] == 59989 && 
b[59990] == 59990 && 
b[59991] == 59991 && 
b[59992] == 59992 && 
b[59993] == 59993 && 
b[59994] == 59994 && 
b[59995] == 59995 && 
b[59996] == 59996 && 
b[59997] == 59997 && 
b[59998] == 59998 && 
b[59999] == 59999 && 
b[60000] == 60000 && 
b[60001] == 60001 && 
b[60002] == 60002 && 
b[60003] == 60003 && 
b[60004] == 60004 && 
b[60005] == 60005 && 
b[60006] == 60006 && 
b[60007] == 60007 && 
b[60008] == 60008 && 
b[60009] == 60009 && 
b[60010] == 60010 && 
b[60011] == 60011 && 
b[60012] == 60012 && 
b[60013] == 60013 && 
b[60014] == 60014 && 
b[60015] == 60015 && 
b[60016] == 60016 && 
b[60017] == 60017 && 
b[60018] == 60018 && 
b[60019] == 60019 && 
b[60020] == 60020 && 
b[60021] == 60021 && 
b[60022] == 60022 && 
b[60023] == 60023 && 
b[60024] == 60024 && 
b[60025] == 60025 && 
b[60026] == 60026 && 
b[60027] == 60027 && 
b[60028] == 60028 && 
b[60029] == 60029 && 
b[60030] == 60030 && 
b[60031] == 60031 && 
b[60032] == 60032 && 
b[60033] == 60033 && 
b[60034] == 60034 && 
b[60035] == 60035 && 
b[60036] == 60036 && 
b[60037] == 60037 && 
b[60038] == 60038 && 
b[60039] == 60039 && 
b[60040] == 60040 && 
b[60041] == 60041 && 
b[60042] == 60042 && 
b[60043] == 60043 && 
b[60044] == 60044 && 
b[60045] == 60045 && 
b[60046] == 60046 && 
b[60047] == 60047 && 
b[60048] == 60048 && 
b[60049] == 60049 && 
b[60050] == 60050 && 
b[60051] == 60051 && 
b[60052] == 60052 && 
b[60053] == 60053 && 
b[60054] == 60054 && 
b[60055] == 60055 && 
b[60056] == 60056 && 
b[60057] == 60057 && 
b[60058] == 60058 && 
b[60059] == 60059 && 
b[60060] == 60060 && 
b[60061] == 60061 && 
b[60062] == 60062 && 
b[60063] == 60063 && 
b[60064] == 60064 && 
b[60065] == 60065 && 
b[60066] == 60066 && 
b[60067] == 60067 && 
b[60068] == 60068 && 
b[60069] == 60069 && 
b[60070] == 60070 && 
b[60071] == 60071 && 
b[60072] == 60072 && 
b[60073] == 60073 && 
b[60074] == 60074 && 
b[60075] == 60075 && 
b[60076] == 60076 && 
b[60077] == 60077 && 
b[60078] == 60078 && 
b[60079] == 60079 && 
b[60080] == 60080 && 
b[60081] == 60081 && 
b[60082] == 60082 && 
b[60083] == 60083 && 
b[60084] == 60084 && 
b[60085] == 60085 && 
b[60086] == 60086 && 
b[60087] == 60087 && 
b[60088] == 60088 && 
b[60089] == 60089 && 
b[60090] == 60090 && 
b[60091] == 60091 && 
b[60092] == 60092 && 
b[60093] == 60093 && 
b[60094] == 60094 && 
b[60095] == 60095 && 
b[60096] == 60096 && 
b[60097] == 60097 && 
b[60098] == 60098 && 
b[60099] == 60099 && 
b[60100] == 60100 && 
b[60101] == 60101 && 
b[60102] == 60102 && 
b[60103] == 60103 && 
b[60104] == 60104 && 
b[60105] == 60105 && 
b[60106] == 60106 && 
b[60107] == 60107 && 
b[60108] == 60108 && 
b[60109] == 60109 && 
b[60110] == 60110 && 
b[60111] == 60111 && 
b[60112] == 60112 && 
b[60113] == 60113 && 
b[60114] == 60114 && 
b[60115] == 60115 && 
b[60116] == 60116 && 
b[60117] == 60117 && 
b[60118] == 60118 && 
b[60119] == 60119 && 
b[60120] == 60120 && 
b[60121] == 60121 && 
b[60122] == 60122 && 
b[60123] == 60123 && 
b[60124] == 60124 && 
b[60125] == 60125 && 
b[60126] == 60126 && 
b[60127] == 60127 && 
b[60128] == 60128 && 
b[60129] == 60129 && 
b[60130] == 60130 && 
b[60131] == 60131 && 
b[60132] == 60132 && 
b[60133] == 60133 && 
b[60134] == 60134 && 
b[60135] == 60135 && 
b[60136] == 60136 && 
b[60137] == 60137 && 
b[60138] == 60138 && 
b[60139] == 60139 && 
b[60140] == 60140 && 
b[60141] == 60141 && 
b[60142] == 60142 && 
b[60143] == 60143 && 
b[60144] == 60144 && 
b[60145] == 60145 && 
b[60146] == 60146 && 
b[60147] == 60147 && 
b[60148] == 60148 && 
b[60149] == 60149 && 
b[60150] == 60150 && 
b[60151] == 60151 && 
b[60152] == 60152 && 
b[60153] == 60153 && 
b[60154] == 60154 && 
b[60155] == 60155 && 
b[60156] == 60156 && 
b[60157] == 60157 && 
b[60158] == 60158 && 
b[60159] == 60159 && 
b[60160] == 60160 && 
b[60161] == 60161 && 
b[60162] == 60162 && 
b[60163] == 60163 && 
b[60164] == 60164 && 
b[60165] == 60165 && 
b[60166] == 60166 && 
b[60167] == 60167 && 
b[60168] == 60168 && 
b[60169] == 60169 && 
b[60170] == 60170 && 
b[60171] == 60171 && 
b[60172] == 60172 && 
b[60173] == 60173 && 
b[60174] == 60174 && 
b[60175] == 60175 && 
b[60176] == 60176 && 
b[60177] == 60177 && 
b[60178] == 60178 && 
b[60179] == 60179 && 
b[60180] == 60180 && 
b[60181] == 60181 && 
b[60182] == 60182 && 
b[60183] == 60183 && 
b[60184] == 60184 && 
b[60185] == 60185 && 
b[60186] == 60186 && 
b[60187] == 60187 && 
b[60188] == 60188 && 
b[60189] == 60189 && 
b[60190] == 60190 && 
b[60191] == 60191 && 
b[60192] == 60192 && 
b[60193] == 60193 && 
b[60194] == 60194 && 
b[60195] == 60195 && 
b[60196] == 60196 && 
b[60197] == 60197 && 
b[60198] == 60198 && 
b[60199] == 60199 && 
b[60200] == 60200 && 
b[60201] == 60201 && 
b[60202] == 60202 && 
b[60203] == 60203 && 
b[60204] == 60204 && 
b[60205] == 60205 && 
b[60206] == 60206 && 
b[60207] == 60207 && 
b[60208] == 60208 && 
b[60209] == 60209 && 
b[60210] == 60210 && 
b[60211] == 60211 && 
b[60212] == 60212 && 
b[60213] == 60213 && 
b[60214] == 60214 && 
b[60215] == 60215 && 
b[60216] == 60216 && 
b[60217] == 60217 && 
b[60218] == 60218 && 
b[60219] == 60219 && 
b[60220] == 60220 && 
b[60221] == 60221 && 
b[60222] == 60222 && 
b[60223] == 60223 && 
b[60224] == 60224 && 
b[60225] == 60225 && 
b[60226] == 60226 && 
b[60227] == 60227 && 
b[60228] == 60228 && 
b[60229] == 60229 && 
b[60230] == 60230 && 
b[60231] == 60231 && 
b[60232] == 60232 && 
b[60233] == 60233 && 
b[60234] == 60234 && 
b[60235] == 60235 && 
b[60236] == 60236 && 
b[60237] == 60237 && 
b[60238] == 60238 && 
b[60239] == 60239 && 
b[60240] == 60240 && 
b[60241] == 60241 && 
b[60242] == 60242 && 
b[60243] == 60243 && 
b[60244] == 60244 && 
b[60245] == 60245 && 
b[60246] == 60246 && 
b[60247] == 60247 && 
b[60248] == 60248 && 
b[60249] == 60249 && 
b[60250] == 60250 && 
b[60251] == 60251 && 
b[60252] == 60252 && 
b[60253] == 60253 && 
b[60254] == 60254 && 
b[60255] == 60255 && 
b[60256] == 60256 && 
b[60257] == 60257 && 
b[60258] == 60258 && 
b[60259] == 60259 && 
b[60260] == 60260 && 
b[60261] == 60261 && 
b[60262] == 60262 && 
b[60263] == 60263 && 
b[60264] == 60264 && 
b[60265] == 60265 && 
b[60266] == 60266 && 
b[60267] == 60267 && 
b[60268] == 60268 && 
b[60269] == 60269 && 
b[60270] == 60270 && 
b[60271] == 60271 && 
b[60272] == 60272 && 
b[60273] == 60273 && 
b[60274] == 60274 && 
b[60275] == 60275 && 
b[60276] == 60276 && 
b[60277] == 60277 && 
b[60278] == 60278 && 
b[60279] == 60279 && 
b[60280] == 60280 && 
b[60281] == 60281 && 
b[60282] == 60282 && 
b[60283] == 60283 && 
b[60284] == 60284 && 
b[60285] == 60285 && 
b[60286] == 60286 && 
b[60287] == 60287 && 
b[60288] == 60288 && 
b[60289] == 60289 && 
b[60290] == 60290 && 
b[60291] == 60291 && 
b[60292] == 60292 && 
b[60293] == 60293 && 
b[60294] == 60294 && 
b[60295] == 60295 && 
b[60296] == 60296 && 
b[60297] == 60297 && 
b[60298] == 60298 && 
b[60299] == 60299 && 
b[60300] == 60300 && 
b[60301] == 60301 && 
b[60302] == 60302 && 
b[60303] == 60303 && 
b[60304] == 60304 && 
b[60305] == 60305 && 
b[60306] == 60306 && 
b[60307] == 60307 && 
b[60308] == 60308 && 
b[60309] == 60309 && 
b[60310] == 60310 && 
b[60311] == 60311 && 
b[60312] == 60312 && 
b[60313] == 60313 && 
b[60314] == 60314 && 
b[60315] == 60315 && 
b[60316] == 60316 && 
b[60317] == 60317 && 
b[60318] == 60318 && 
b[60319] == 60319 && 
b[60320] == 60320 && 
b[60321] == 60321 && 
b[60322] == 60322 && 
b[60323] == 60323 && 
b[60324] == 60324 && 
b[60325] == 60325 && 
b[60326] == 60326 && 
b[60327] == 60327 && 
b[60328] == 60328 && 
b[60329] == 60329 && 
b[60330] == 60330 && 
b[60331] == 60331 && 
b[60332] == 60332 && 
b[60333] == 60333 && 
b[60334] == 60334 && 
b[60335] == 60335 && 
b[60336] == 60336 && 
b[60337] == 60337 && 
b[60338] == 60338 && 
b[60339] == 60339 && 
b[60340] == 60340 && 
b[60341] == 60341 && 
b[60342] == 60342 && 
b[60343] == 60343 && 
b[60344] == 60344 && 
b[60345] == 60345 && 
b[60346] == 60346 && 
b[60347] == 60347 && 
b[60348] == 60348 && 
b[60349] == 60349 && 
b[60350] == 60350 && 
b[60351] == 60351 && 
b[60352] == 60352 && 
b[60353] == 60353 && 
b[60354] == 60354 && 
b[60355] == 60355 && 
b[60356] == 60356 && 
b[60357] == 60357 && 
b[60358] == 60358 && 
b[60359] == 60359 && 
b[60360] == 60360 && 
b[60361] == 60361 && 
b[60362] == 60362 && 
b[60363] == 60363 && 
b[60364] == 60364 && 
b[60365] == 60365 && 
b[60366] == 60366 && 
b[60367] == 60367 && 
b[60368] == 60368 && 
b[60369] == 60369 && 
b[60370] == 60370 && 
b[60371] == 60371 && 
b[60372] == 60372 && 
b[60373] == 60373 && 
b[60374] == 60374 && 
b[60375] == 60375 && 
b[60376] == 60376 && 
b[60377] == 60377 && 
b[60378] == 60378 && 
b[60379] == 60379 && 
b[60380] == 60380 && 
b[60381] == 60381 && 
b[60382] == 60382 && 
b[60383] == 60383 && 
b[60384] == 60384 && 
b[60385] == 60385 && 
b[60386] == 60386 && 
b[60387] == 60387 && 
b[60388] == 60388 && 
b[60389] == 60389 && 
b[60390] == 60390 && 
b[60391] == 60391 && 
b[60392] == 60392 && 
b[60393] == 60393 && 
b[60394] == 60394 && 
b[60395] == 60395 && 
b[60396] == 60396 && 
b[60397] == 60397 && 
b[60398] == 60398 && 
b[60399] == 60399 && 
b[60400] == 60400 && 
b[60401] == 60401 && 
b[60402] == 60402 && 
b[60403] == 60403 && 
b[60404] == 60404 && 
b[60405] == 60405 && 
b[60406] == 60406 && 
b[60407] == 60407 && 
b[60408] == 60408 && 
b[60409] == 60409 && 
b[60410] == 60410 && 
b[60411] == 60411 && 
b[60412] == 60412 && 
b[60413] == 60413 && 
b[60414] == 60414 && 
b[60415] == 60415 && 
b[60416] == 60416 && 
b[60417] == 60417 && 
b[60418] == 60418 && 
b[60419] == 60419 && 
b[60420] == 60420 && 
b[60421] == 60421 && 
b[60422] == 60422 && 
b[60423] == 60423 && 
b[60424] == 60424 && 
b[60425] == 60425 && 
b[60426] == 60426 && 
b[60427] == 60427 && 
b[60428] == 60428 && 
b[60429] == 60429 && 
b[60430] == 60430 && 
b[60431] == 60431 && 
b[60432] == 60432 && 
b[60433] == 60433 && 
b[60434] == 60434 && 
b[60435] == 60435 && 
b[60436] == 60436 && 
b[60437] == 60437 && 
b[60438] == 60438 && 
b[60439] == 60439 && 
b[60440] == 60440 && 
b[60441] == 60441 && 
b[60442] == 60442 && 
b[60443] == 60443 && 
b[60444] == 60444 && 
b[60445] == 60445 && 
b[60446] == 60446 && 
b[60447] == 60447 && 
b[60448] == 60448 && 
b[60449] == 60449 && 
b[60450] == 60450 && 
b[60451] == 60451 && 
b[60452] == 60452 && 
b[60453] == 60453 && 
b[60454] == 60454 && 
b[60455] == 60455 && 
b[60456] == 60456 && 
b[60457] == 60457 && 
b[60458] == 60458 && 
b[60459] == 60459 && 
b[60460] == 60460 && 
b[60461] == 60461 && 
b[60462] == 60462 && 
b[60463] == 60463 && 
b[60464] == 60464 && 
b[60465] == 60465 && 
b[60466] == 60466 && 
b[60467] == 60467 && 
b[60468] == 60468 && 
b[60469] == 60469 && 
b[60470] == 60470 && 
b[60471] == 60471 && 
b[60472] == 60472 && 
b[60473] == 60473 && 
b[60474] == 60474 && 
b[60475] == 60475 && 
b[60476] == 60476 && 
b[60477] == 60477 && 
b[60478] == 60478 && 
b[60479] == 60479 && 
b[60480] == 60480 && 
b[60481] == 60481 && 
b[60482] == 60482 && 
b[60483] == 60483 && 
b[60484] == 60484 && 
b[60485] == 60485 && 
b[60486] == 60486 && 
b[60487] == 60487 && 
b[60488] == 60488 && 
b[60489] == 60489 && 
b[60490] == 60490 && 
b[60491] == 60491 && 
b[60492] == 60492 && 
b[60493] == 60493 && 
b[60494] == 60494 && 
b[60495] == 60495 && 
b[60496] == 60496 && 
b[60497] == 60497 && 
b[60498] == 60498 && 
b[60499] == 60499 && 
b[60500] == 60500 && 
b[60501] == 60501 && 
b[60502] == 60502 && 
b[60503] == 60503 && 
b[60504] == 60504 && 
b[60505] == 60505 && 
b[60506] == 60506 && 
b[60507] == 60507 && 
b[60508] == 60508 && 
b[60509] == 60509 && 
b[60510] == 60510 && 
b[60511] == 60511 && 
b[60512] == 60512 && 
b[60513] == 60513 && 
b[60514] == 60514 && 
b[60515] == 60515 && 
b[60516] == 60516 && 
b[60517] == 60517 && 
b[60518] == 60518 && 
b[60519] == 60519 && 
b[60520] == 60520 && 
b[60521] == 60521 && 
b[60522] == 60522 && 
b[60523] == 60523 && 
b[60524] == 60524 && 
b[60525] == 60525 && 
b[60526] == 60526 && 
b[60527] == 60527 && 
b[60528] == 60528 && 
b[60529] == 60529 && 
b[60530] == 60530 && 
b[60531] == 60531 && 
b[60532] == 60532 && 
b[60533] == 60533 && 
b[60534] == 60534 && 
b[60535] == 60535 && 
b[60536] == 60536 && 
b[60537] == 60537 && 
b[60538] == 60538 && 
b[60539] == 60539 && 
b[60540] == 60540 && 
b[60541] == 60541 && 
b[60542] == 60542 && 
b[60543] == 60543 && 
b[60544] == 60544 && 
b[60545] == 60545 && 
b[60546] == 60546 && 
b[60547] == 60547 && 
b[60548] == 60548 && 
b[60549] == 60549 && 
b[60550] == 60550 && 
b[60551] == 60551 && 
b[60552] == 60552 && 
b[60553] == 60553 && 
b[60554] == 60554 && 
b[60555] == 60555 && 
b[60556] == 60556 && 
b[60557] == 60557 && 
b[60558] == 60558 && 
b[60559] == 60559 && 
b[60560] == 60560 && 
b[60561] == 60561 && 
b[60562] == 60562 && 
b[60563] == 60563 && 
b[60564] == 60564 && 
b[60565] == 60565 && 
b[60566] == 60566 && 
b[60567] == 60567 && 
b[60568] == 60568 && 
b[60569] == 60569 && 
b[60570] == 60570 && 
b[60571] == 60571 && 
b[60572] == 60572 && 
b[60573] == 60573 && 
b[60574] == 60574 && 
b[60575] == 60575 && 
b[60576] == 60576 && 
b[60577] == 60577 && 
b[60578] == 60578 && 
b[60579] == 60579 && 
b[60580] == 60580 && 
b[60581] == 60581 && 
b[60582] == 60582 && 
b[60583] == 60583 && 
b[60584] == 60584 && 
b[60585] == 60585 && 
b[60586] == 60586 && 
b[60587] == 60587 && 
b[60588] == 60588 && 
b[60589] == 60589 && 
b[60590] == 60590 && 
b[60591] == 60591 && 
b[60592] == 60592 && 
b[60593] == 60593 && 
b[60594] == 60594 && 
b[60595] == 60595 && 
b[60596] == 60596 && 
b[60597] == 60597 && 
b[60598] == 60598 && 
b[60599] == 60599 && 
b[60600] == 60600 && 
b[60601] == 60601 && 
b[60602] == 60602 && 
b[60603] == 60603 && 
b[60604] == 60604 && 
b[60605] == 60605 && 
b[60606] == 60606 && 
b[60607] == 60607 && 
b[60608] == 60608 && 
b[60609] == 60609 && 
b[60610] == 60610 && 
b[60611] == 60611 && 
b[60612] == 60612 && 
b[60613] == 60613 && 
b[60614] == 60614 && 
b[60615] == 60615 && 
b[60616] == 60616 && 
b[60617] == 60617 && 
b[60618] == 60618 && 
b[60619] == 60619 && 
b[60620] == 60620 && 
b[60621] == 60621 && 
b[60622] == 60622 && 
b[60623] == 60623 && 
b[60624] == 60624 && 
b[60625] == 60625 && 
b[60626] == 60626 && 
b[60627] == 60627 && 
b[60628] == 60628 && 
b[60629] == 60629 && 
b[60630] == 60630 && 
b[60631] == 60631 && 
b[60632] == 60632 && 
b[60633] == 60633 && 
b[60634] == 60634 && 
b[60635] == 60635 && 
b[60636] == 60636 && 
b[60637] == 60637 && 
b[60638] == 60638 && 
b[60639] == 60639 && 
b[60640] == 60640 && 
b[60641] == 60641 && 
b[60642] == 60642 && 
b[60643] == 60643 && 
b[60644] == 60644 && 
b[60645] == 60645 && 
b[60646] == 60646 && 
b[60647] == 60647 && 
b[60648] == 60648 && 
b[60649] == 60649 && 
b[60650] == 60650 && 
b[60651] == 60651 && 
b[60652] == 60652 && 
b[60653] == 60653 && 
b[60654] == 60654 && 
b[60655] == 60655 && 
b[60656] == 60656 && 
b[60657] == 60657 && 
b[60658] == 60658 && 
b[60659] == 60659 && 
b[60660] == 60660 && 
b[60661] == 60661 && 
b[60662] == 60662 && 
b[60663] == 60663 && 
b[60664] == 60664 && 
b[60665] == 60665 && 
b[60666] == 60666 && 
b[60667] == 60667 && 
b[60668] == 60668 && 
b[60669] == 60669 && 
b[60670] == 60670 && 
b[60671] == 60671 && 
b[60672] == 60672 && 
b[60673] == 60673 && 
b[60674] == 60674 && 
b[60675] == 60675 && 
b[60676] == 60676 && 
b[60677] == 60677 && 
b[60678] == 60678 && 
b[60679] == 60679 && 
b[60680] == 60680 && 
b[60681] == 60681 && 
b[60682] == 60682 && 
b[60683] == 60683 && 
b[60684] == 60684 && 
b[60685] == 60685 && 
b[60686] == 60686 && 
b[60687] == 60687 && 
b[60688] == 60688 && 
b[60689] == 60689 && 
b[60690] == 60690 && 
b[60691] == 60691 && 
b[60692] == 60692 && 
b[60693] == 60693 && 
b[60694] == 60694 && 
b[60695] == 60695 && 
b[60696] == 60696 && 
b[60697] == 60697 && 
b[60698] == 60698 && 
b[60699] == 60699 && 
b[60700] == 60700 && 
b[60701] == 60701 && 
b[60702] == 60702 && 
b[60703] == 60703 && 
b[60704] == 60704 && 
b[60705] == 60705 && 
b[60706] == 60706 && 
b[60707] == 60707 && 
b[60708] == 60708 && 
b[60709] == 60709 && 
b[60710] == 60710 && 
b[60711] == 60711 && 
b[60712] == 60712 && 
b[60713] == 60713 && 
b[60714] == 60714 && 
b[60715] == 60715 && 
b[60716] == 60716 && 
b[60717] == 60717 && 
b[60718] == 60718 && 
b[60719] == 60719 && 
b[60720] == 60720 && 
b[60721] == 60721 && 
b[60722] == 60722 && 
b[60723] == 60723 && 
b[60724] == 60724 && 
b[60725] == 60725 && 
b[60726] == 60726 && 
b[60727] == 60727 && 
b[60728] == 60728 && 
b[60729] == 60729 && 
b[60730] == 60730 && 
b[60731] == 60731 && 
b[60732] == 60732 && 
b[60733] == 60733 && 
b[60734] == 60734 && 
b[60735] == 60735 && 
b[60736] == 60736 && 
b[60737] == 60737 && 
b[60738] == 60738 && 
b[60739] == 60739 && 
b[60740] == 60740 && 
b[60741] == 60741 && 
b[60742] == 60742 && 
b[60743] == 60743 && 
b[60744] == 60744 && 
b[60745] == 60745 && 
b[60746] == 60746 && 
b[60747] == 60747 && 
b[60748] == 60748 && 
b[60749] == 60749 && 
b[60750] == 60750 && 
b[60751] == 60751 && 
b[60752] == 60752 && 
b[60753] == 60753 && 
b[60754] == 60754 && 
b[60755] == 60755 && 
b[60756] == 60756 && 
b[60757] == 60757 && 
b[60758] == 60758 && 
b[60759] == 60759 && 
b[60760] == 60760 && 
b[60761] == 60761 && 
b[60762] == 60762 && 
b[60763] == 60763 && 
b[60764] == 60764 && 
b[60765] == 60765 && 
b[60766] == 60766 && 
b[60767] == 60767 && 
b[60768] == 60768 && 
b[60769] == 60769 && 
b[60770] == 60770 && 
b[60771] == 60771 && 
b[60772] == 60772 && 
b[60773] == 60773 && 
b[60774] == 60774 && 
b[60775] == 60775 && 
b[60776] == 60776 && 
b[60777] == 60777 && 
b[60778] == 60778 && 
b[60779] == 60779 && 
b[60780] == 60780 && 
b[60781] == 60781 && 
b[60782] == 60782 && 
b[60783] == 60783 && 
b[60784] == 60784 && 
b[60785] == 60785 && 
b[60786] == 60786 && 
b[60787] == 60787 && 
b[60788] == 60788 && 
b[60789] == 60789 && 
b[60790] == 60790 && 
b[60791] == 60791 && 
b[60792] == 60792 && 
b[60793] == 60793 && 
b[60794] == 60794 && 
b[60795] == 60795 && 
b[60796] == 60796 && 
b[60797] == 60797 && 
b[60798] == 60798 && 
b[60799] == 60799 && 
b[60800] == 60800 && 
b[60801] == 60801 && 
b[60802] == 60802 && 
b[60803] == 60803 && 
b[60804] == 60804 && 
b[60805] == 60805 && 
b[60806] == 60806 && 
b[60807] == 60807 && 
b[60808] == 60808 && 
b[60809] == 60809 && 
b[60810] == 60810 && 
b[60811] == 60811 && 
b[60812] == 60812 && 
b[60813] == 60813 && 
b[60814] == 60814 && 
b[60815] == 60815 && 
b[60816] == 60816 && 
b[60817] == 60817 && 
b[60818] == 60818 && 
b[60819] == 60819 && 
b[60820] == 60820 && 
b[60821] == 60821 && 
b[60822] == 60822 && 
b[60823] == 60823 && 
b[60824] == 60824 && 
b[60825] == 60825 && 
b[60826] == 60826 && 
b[60827] == 60827 && 
b[60828] == 60828 && 
b[60829] == 60829 && 
b[60830] == 60830 && 
b[60831] == 60831 && 
b[60832] == 60832 && 
b[60833] == 60833 && 
b[60834] == 60834 && 
b[60835] == 60835 && 
b[60836] == 60836 && 
b[60837] == 60837 && 
b[60838] == 60838 && 
b[60839] == 60839 && 
b[60840] == 60840 && 
b[60841] == 60841 && 
b[60842] == 60842 && 
b[60843] == 60843 && 
b[60844] == 60844 && 
b[60845] == 60845 && 
b[60846] == 60846 && 
b[60847] == 60847 && 
b[60848] == 60848 && 
b[60849] == 60849 && 
b[60850] == 60850 && 
b[60851] == 60851 && 
b[60852] == 60852 && 
b[60853] == 60853 && 
b[60854] == 60854 && 
b[60855] == 60855 && 
b[60856] == 60856 && 
b[60857] == 60857 && 
b[60858] == 60858 && 
b[60859] == 60859 && 
b[60860] == 60860 && 
b[60861] == 60861 && 
b[60862] == 60862 && 
b[60863] == 60863 && 
b[60864] == 60864 && 
b[60865] == 60865 && 
b[60866] == 60866 && 
b[60867] == 60867 && 
b[60868] == 60868 && 
b[60869] == 60869 && 
b[60870] == 60870 && 
b[60871] == 60871 && 
b[60872] == 60872 && 
b[60873] == 60873 && 
b[60874] == 60874 && 
b[60875] == 60875 && 
b[60876] == 60876 && 
b[60877] == 60877 && 
b[60878] == 60878 && 
b[60879] == 60879 && 
b[60880] == 60880 && 
b[60881] == 60881 && 
b[60882] == 60882 && 
b[60883] == 60883 && 
b[60884] == 60884 && 
b[60885] == 60885 && 
b[60886] == 60886 && 
b[60887] == 60887 && 
b[60888] == 60888 && 
b[60889] == 60889 && 
b[60890] == 60890 && 
b[60891] == 60891 && 
b[60892] == 60892 && 
b[60893] == 60893 && 
b[60894] == 60894 && 
b[60895] == 60895 && 
b[60896] == 60896 && 
b[60897] == 60897 && 
b[60898] == 60898 && 
b[60899] == 60899 && 
b[60900] == 60900 && 
b[60901] == 60901 && 
b[60902] == 60902 && 
b[60903] == 60903 && 
b[60904] == 60904 && 
b[60905] == 60905 && 
b[60906] == 60906 && 
b[60907] == 60907 && 
b[60908] == 60908 && 
b[60909] == 60909 && 
b[60910] == 60910 && 
b[60911] == 60911 && 
b[60912] == 60912 && 
b[60913] == 60913 && 
b[60914] == 60914 && 
b[60915] == 60915 && 
b[60916] == 60916 && 
b[60917] == 60917 && 
b[60918] == 60918 && 
b[60919] == 60919 && 
b[60920] == 60920 && 
b[60921] == 60921 && 
b[60922] == 60922 && 
b[60923] == 60923 && 
b[60924] == 60924 && 
b[60925] == 60925 && 
b[60926] == 60926 && 
b[60927] == 60927 && 
b[60928] == 60928 && 
b[60929] == 60929 && 
b[60930] == 60930 && 
b[60931] == 60931 && 
b[60932] == 60932 && 
b[60933] == 60933 && 
b[60934] == 60934 && 
b[60935] == 60935 && 
b[60936] == 60936 && 
b[60937] == 60937 && 
b[60938] == 60938 && 
b[60939] == 60939 && 
b[60940] == 60940 && 
b[60941] == 60941 && 
b[60942] == 60942 && 
b[60943] == 60943 && 
b[60944] == 60944 && 
b[60945] == 60945 && 
b[60946] == 60946 && 
b[60947] == 60947 && 
b[60948] == 60948 && 
b[60949] == 60949 && 
b[60950] == 60950 && 
b[60951] == 60951 && 
b[60952] == 60952 && 
b[60953] == 60953 && 
b[60954] == 60954 && 
b[60955] == 60955 && 
b[60956] == 60956 && 
b[60957] == 60957 && 
b[60958] == 60958 && 
b[60959] == 60959 && 
b[60960] == 60960 && 
b[60961] == 60961 && 
b[60962] == 60962 && 
b[60963] == 60963 && 
b[60964] == 60964 && 
b[60965] == 60965 && 
b[60966] == 60966 && 
b[60967] == 60967 && 
b[60968] == 60968 && 
b[60969] == 60969 && 
b[60970] == 60970 && 
b[60971] == 60971 && 
b[60972] == 60972 && 
b[60973] == 60973 && 
b[60974] == 60974 && 
b[60975] == 60975 && 
b[60976] == 60976 && 
b[60977] == 60977 && 
b[60978] == 60978 && 
b[60979] == 60979 && 
b[60980] == 60980 && 
b[60981] == 60981 && 
b[60982] == 60982 && 
b[60983] == 60983 && 
b[60984] == 60984 && 
b[60985] == 60985 && 
b[60986] == 60986 && 
b[60987] == 60987 && 
b[60988] == 60988 && 
b[60989] == 60989 && 
b[60990] == 60990 && 
b[60991] == 60991 && 
b[60992] == 60992 && 
b[60993] == 60993 && 
b[60994] == 60994 && 
b[60995] == 60995 && 
b[60996] == 60996 && 
b[60997] == 60997 && 
b[60998] == 60998 && 
b[60999] == 60999 && 
b[61000] == 61000 && 
b[61001] == 61001 && 
b[61002] == 61002 && 
b[61003] == 61003 && 
b[61004] == 61004 && 
b[61005] == 61005 && 
b[61006] == 61006 && 
b[61007] == 61007 && 
b[61008] == 61008 && 
b[61009] == 61009 && 
b[61010] == 61010 && 
b[61011] == 61011 && 
b[61012] == 61012 && 
b[61013] == 61013 && 
b[61014] == 61014 && 
b[61015] == 61015 && 
b[61016] == 61016 && 
b[61017] == 61017 && 
b[61018] == 61018 && 
b[61019] == 61019 && 
b[61020] == 61020 && 
b[61021] == 61021 && 
b[61022] == 61022 && 
b[61023] == 61023 && 
b[61024] == 61024 && 
b[61025] == 61025 && 
b[61026] == 61026 && 
b[61027] == 61027 && 
b[61028] == 61028 && 
b[61029] == 61029 && 
b[61030] == 61030 && 
b[61031] == 61031 && 
b[61032] == 61032 && 
b[61033] == 61033 && 
b[61034] == 61034 && 
b[61035] == 61035 && 
b[61036] == 61036 && 
b[61037] == 61037 && 
b[61038] == 61038 && 
b[61039] == 61039 && 
b[61040] == 61040 && 
b[61041] == 61041 && 
b[61042] == 61042 && 
b[61043] == 61043 && 
b[61044] == 61044 && 
b[61045] == 61045 && 
b[61046] == 61046 && 
b[61047] == 61047 && 
b[61048] == 61048 && 
b[61049] == 61049 && 
b[61050] == 61050 && 
b[61051] == 61051 && 
b[61052] == 61052 && 
b[61053] == 61053 && 
b[61054] == 61054 && 
b[61055] == 61055 && 
b[61056] == 61056 && 
b[61057] == 61057 && 
b[61058] == 61058 && 
b[61059] == 61059 && 
b[61060] == 61060 && 
b[61061] == 61061 && 
b[61062] == 61062 && 
b[61063] == 61063 && 
b[61064] == 61064 && 
b[61065] == 61065 && 
b[61066] == 61066 && 
b[61067] == 61067 && 
b[61068] == 61068 && 
b[61069] == 61069 && 
b[61070] == 61070 && 
b[61071] == 61071 && 
b[61072] == 61072 && 
b[61073] == 61073 && 
b[61074] == 61074 && 
b[61075] == 61075 && 
b[61076] == 61076 && 
b[61077] == 61077 && 
b[61078] == 61078 && 
b[61079] == 61079 && 
b[61080] == 61080 && 
b[61081] == 61081 && 
b[61082] == 61082 && 
b[61083] == 61083 && 
b[61084] == 61084 && 
b[61085] == 61085 && 
b[61086] == 61086 && 
b[61087] == 61087 && 
b[61088] == 61088 && 
b[61089] == 61089 && 
b[61090] == 61090 && 
b[61091] == 61091 && 
b[61092] == 61092 && 
b[61093] == 61093 && 
b[61094] == 61094 && 
b[61095] == 61095 && 
b[61096] == 61096 && 
b[61097] == 61097 && 
b[61098] == 61098 && 
b[61099] == 61099 && 
b[61100] == 61100 && 
b[61101] == 61101 && 
b[61102] == 61102 && 
b[61103] == 61103 && 
b[61104] == 61104 && 
b[61105] == 61105 && 
b[61106] == 61106 && 
b[61107] == 61107 && 
b[61108] == 61108 && 
b[61109] == 61109 && 
b[61110] == 61110 && 
b[61111] == 61111 && 
b[61112] == 61112 && 
b[61113] == 61113 && 
b[61114] == 61114 && 
b[61115] == 61115 && 
b[61116] == 61116 && 
b[61117] == 61117 && 
b[61118] == 61118 && 
b[61119] == 61119 && 
b[61120] == 61120 && 
b[61121] == 61121 && 
b[61122] == 61122 && 
b[61123] == 61123 && 
b[61124] == 61124 && 
b[61125] == 61125 && 
b[61126] == 61126 && 
b[61127] == 61127 && 
b[61128] == 61128 && 
b[61129] == 61129 && 
b[61130] == 61130 && 
b[61131] == 61131 && 
b[61132] == 61132 && 
b[61133] == 61133 && 
b[61134] == 61134 && 
b[61135] == 61135 && 
b[61136] == 61136 && 
b[61137] == 61137 && 
b[61138] == 61138 && 
b[61139] == 61139 && 
b[61140] == 61140 && 
b[61141] == 61141 && 
b[61142] == 61142 && 
b[61143] == 61143 && 
b[61144] == 61144 && 
b[61145] == 61145 && 
b[61146] == 61146 && 
b[61147] == 61147 && 
b[61148] == 61148 && 
b[61149] == 61149 && 
b[61150] == 61150 && 
b[61151] == 61151 && 
b[61152] == 61152 && 
b[61153] == 61153 && 
b[61154] == 61154 && 
b[61155] == 61155 && 
b[61156] == 61156 && 
b[61157] == 61157 && 
b[61158] == 61158 && 
b[61159] == 61159 && 
b[61160] == 61160 && 
b[61161] == 61161 && 
b[61162] == 61162 && 
b[61163] == 61163 && 
b[61164] == 61164 && 
b[61165] == 61165 && 
b[61166] == 61166 && 
b[61167] == 61167 && 
b[61168] == 61168 && 
b[61169] == 61169 && 
b[61170] == 61170 && 
b[61171] == 61171 && 
b[61172] == 61172 && 
b[61173] == 61173 && 
b[61174] == 61174 && 
b[61175] == 61175 && 
b[61176] == 61176 && 
b[61177] == 61177 && 
b[61178] == 61178 && 
b[61179] == 61179 && 
b[61180] == 61180 && 
b[61181] == 61181 && 
b[61182] == 61182 && 
b[61183] == 61183 && 
b[61184] == 61184 && 
b[61185] == 61185 && 
b[61186] == 61186 && 
b[61187] == 61187 && 
b[61188] == 61188 && 
b[61189] == 61189 && 
b[61190] == 61190 && 
b[61191] == 61191 && 
b[61192] == 61192 && 
b[61193] == 61193 && 
b[61194] == 61194 && 
b[61195] == 61195 && 
b[61196] == 61196 && 
b[61197] == 61197 && 
b[61198] == 61198 && 
b[61199] == 61199 && 
b[61200] == 61200 && 
b[61201] == 61201 && 
b[61202] == 61202 && 
b[61203] == 61203 && 
b[61204] == 61204 && 
b[61205] == 61205 && 
b[61206] == 61206 && 
b[61207] == 61207 && 
b[61208] == 61208 && 
b[61209] == 61209 && 
b[61210] == 61210 && 
b[61211] == 61211 && 
b[61212] == 61212 && 
b[61213] == 61213 && 
b[61214] == 61214 && 
b[61215] == 61215 && 
b[61216] == 61216 && 
b[61217] == 61217 && 
b[61218] == 61218 && 
b[61219] == 61219 && 
b[61220] == 61220 && 
b[61221] == 61221 && 
b[61222] == 61222 && 
b[61223] == 61223 && 
b[61224] == 61224 && 
b[61225] == 61225 && 
b[61226] == 61226 && 
b[61227] == 61227 && 
b[61228] == 61228 && 
b[61229] == 61229 && 
b[61230] == 61230 && 
b[61231] == 61231 && 
b[61232] == 61232 && 
b[61233] == 61233 && 
b[61234] == 61234 && 
b[61235] == 61235 && 
b[61236] == 61236 && 
b[61237] == 61237 && 
b[61238] == 61238 && 
b[61239] == 61239 && 
b[61240] == 61240 && 
b[61241] == 61241 && 
b[61242] == 61242 && 
b[61243] == 61243 && 
b[61244] == 61244 && 
b[61245] == 61245 && 
b[61246] == 61246 && 
b[61247] == 61247 && 
b[61248] == 61248 && 
b[61249] == 61249 && 
b[61250] == 61250 && 
b[61251] == 61251 && 
b[61252] == 61252 && 
b[61253] == 61253 && 
b[61254] == 61254 && 
b[61255] == 61255 && 
b[61256] == 61256 && 
b[61257] == 61257 && 
b[61258] == 61258 && 
b[61259] == 61259 && 
b[61260] == 61260 && 
b[61261] == 61261 && 
b[61262] == 61262 && 
b[61263] == 61263 && 
b[61264] == 61264 && 
b[61265] == 61265 && 
b[61266] == 61266 && 
b[61267] == 61267 && 
b[61268] == 61268 && 
b[61269] == 61269 && 
b[61270] == 61270 && 
b[61271] == 61271 && 
b[61272] == 61272 && 
b[61273] == 61273 && 
b[61274] == 61274 && 
b[61275] == 61275 && 
b[61276] == 61276 && 
b[61277] == 61277 && 
b[61278] == 61278 && 
b[61279] == 61279 && 
b[61280] == 61280 && 
b[61281] == 61281 && 
b[61282] == 61282 && 
b[61283] == 61283 && 
b[61284] == 61284 && 
b[61285] == 61285 && 
b[61286] == 61286 && 
b[61287] == 61287 && 
b[61288] == 61288 && 
b[61289] == 61289 && 
b[61290] == 61290 && 
b[61291] == 61291 && 
b[61292] == 61292 && 
b[61293] == 61293 && 
b[61294] == 61294 && 
b[61295] == 61295 && 
b[61296] == 61296 && 
b[61297] == 61297 && 
b[61298] == 61298 && 
b[61299] == 61299 && 
b[61300] == 61300 && 
b[61301] == 61301 && 
b[61302] == 61302 && 
b[61303] == 61303 && 
b[61304] == 61304 && 
b[61305] == 61305 && 
b[61306] == 61306 && 
b[61307] == 61307 && 
b[61308] == 61308 && 
b[61309] == 61309 && 
b[61310] == 61310 && 
b[61311] == 61311 && 
b[61312] == 61312 && 
b[61313] == 61313 && 
b[61314] == 61314 && 
b[61315] == 61315 && 
b[61316] == 61316 && 
b[61317] == 61317 && 
b[61318] == 61318 && 
b[61319] == 61319 && 
b[61320] == 61320 && 
b[61321] == 61321 && 
b[61322] == 61322 && 
b[61323] == 61323 && 
b[61324] == 61324 && 
b[61325] == 61325 && 
b[61326] == 61326 && 
b[61327] == 61327 && 
b[61328] == 61328 && 
b[61329] == 61329 && 
b[61330] == 61330 && 
b[61331] == 61331 && 
b[61332] == 61332 && 
b[61333] == 61333 && 
b[61334] == 61334 && 
b[61335] == 61335 && 
b[61336] == 61336 && 
b[61337] == 61337 && 
b[61338] == 61338 && 
b[61339] == 61339 && 
b[61340] == 61340 && 
b[61341] == 61341 && 
b[61342] == 61342 && 
b[61343] == 61343 && 
b[61344] == 61344 && 
b[61345] == 61345 && 
b[61346] == 61346 && 
b[61347] == 61347 && 
b[61348] == 61348 && 
b[61349] == 61349 && 
b[61350] == 61350 && 
b[61351] == 61351 && 
b[61352] == 61352 && 
b[61353] == 61353 && 
b[61354] == 61354 && 
b[61355] == 61355 && 
b[61356] == 61356 && 
b[61357] == 61357 && 
b[61358] == 61358 && 
b[61359] == 61359 && 
b[61360] == 61360 && 
b[61361] == 61361 && 
b[61362] == 61362 && 
b[61363] == 61363 && 
b[61364] == 61364 && 
b[61365] == 61365 && 
b[61366] == 61366 && 
b[61367] == 61367 && 
b[61368] == 61368 && 
b[61369] == 61369 && 
b[61370] == 61370 && 
b[61371] == 61371 && 
b[61372] == 61372 && 
b[61373] == 61373 && 
b[61374] == 61374 && 
b[61375] == 61375 && 
b[61376] == 61376 && 
b[61377] == 61377 && 
b[61378] == 61378 && 
b[61379] == 61379 && 
b[61380] == 61380 && 
b[61381] == 61381 && 
b[61382] == 61382 && 
b[61383] == 61383 && 
b[61384] == 61384 && 
b[61385] == 61385 && 
b[61386] == 61386 && 
b[61387] == 61387 && 
b[61388] == 61388 && 
b[61389] == 61389 && 
b[61390] == 61390 && 
b[61391] == 61391 && 
b[61392] == 61392 && 
b[61393] == 61393 && 
b[61394] == 61394 && 
b[61395] == 61395 && 
b[61396] == 61396 && 
b[61397] == 61397 && 
b[61398] == 61398 && 
b[61399] == 61399 && 
b[61400] == 61400 && 
b[61401] == 61401 && 
b[61402] == 61402 && 
b[61403] == 61403 && 
b[61404] == 61404 && 
b[61405] == 61405 && 
b[61406] == 61406 && 
b[61407] == 61407 && 
b[61408] == 61408 && 
b[61409] == 61409 && 
b[61410] == 61410 && 
b[61411] == 61411 && 
b[61412] == 61412 && 
b[61413] == 61413 && 
b[61414] == 61414 && 
b[61415] == 61415 && 
b[61416] == 61416 && 
b[61417] == 61417 && 
b[61418] == 61418 && 
b[61419] == 61419 && 
b[61420] == 61420 && 
b[61421] == 61421 && 
b[61422] == 61422 && 
b[61423] == 61423 && 
b[61424] == 61424 && 
b[61425] == 61425 && 
b[61426] == 61426 && 
b[61427] == 61427 && 
b[61428] == 61428 && 
b[61429] == 61429 && 
b[61430] == 61430 && 
b[61431] == 61431 && 
b[61432] == 61432 && 
b[61433] == 61433 && 
b[61434] == 61434 && 
b[61435] == 61435 && 
b[61436] == 61436 && 
b[61437] == 61437 && 
b[61438] == 61438 && 
b[61439] == 61439 && 
b[61440] == 61440 && 
b[61441] == 61441 && 
b[61442] == 61442 && 
b[61443] == 61443 && 
b[61444] == 61444 && 
b[61445] == 61445 && 
b[61446] == 61446 && 
b[61447] == 61447 && 
b[61448] == 61448 && 
b[61449] == 61449 && 
b[61450] == 61450 && 
b[61451] == 61451 && 
b[61452] == 61452 && 
b[61453] == 61453 && 
b[61454] == 61454 && 
b[61455] == 61455 && 
b[61456] == 61456 && 
b[61457] == 61457 && 
b[61458] == 61458 && 
b[61459] == 61459 && 
b[61460] == 61460 && 
b[61461] == 61461 && 
b[61462] == 61462 && 
b[61463] == 61463 && 
b[61464] == 61464 && 
b[61465] == 61465 && 
b[61466] == 61466 && 
b[61467] == 61467 && 
b[61468] == 61468 && 
b[61469] == 61469 && 
b[61470] == 61470 && 
b[61471] == 61471 && 
b[61472] == 61472 && 
b[61473] == 61473 && 
b[61474] == 61474 && 
b[61475] == 61475 && 
b[61476] == 61476 && 
b[61477] == 61477 && 
b[61478] == 61478 && 
b[61479] == 61479 && 
b[61480] == 61480 && 
b[61481] == 61481 && 
b[61482] == 61482 && 
b[61483] == 61483 && 
b[61484] == 61484 && 
b[61485] == 61485 && 
b[61486] == 61486 && 
b[61487] == 61487 && 
b[61488] == 61488 && 
b[61489] == 61489 && 
b[61490] == 61490 && 
b[61491] == 61491 && 
b[61492] == 61492 && 
b[61493] == 61493 && 
b[61494] == 61494 && 
b[61495] == 61495 && 
b[61496] == 61496 && 
b[61497] == 61497 && 
b[61498] == 61498 && 
b[61499] == 61499 && 
b[61500] == 61500 && 
b[61501] == 61501 && 
b[61502] == 61502 && 
b[61503] == 61503 && 
b[61504] == 61504 && 
b[61505] == 61505 && 
b[61506] == 61506 && 
b[61507] == 61507 && 
b[61508] == 61508 && 
b[61509] == 61509 && 
b[61510] == 61510 && 
b[61511] == 61511 && 
b[61512] == 61512 && 
b[61513] == 61513 && 
b[61514] == 61514 && 
b[61515] == 61515 && 
b[61516] == 61516 && 
b[61517] == 61517 && 
b[61518] == 61518 && 
b[61519] == 61519 && 
b[61520] == 61520 && 
b[61521] == 61521 && 
b[61522] == 61522 && 
b[61523] == 61523 && 
b[61524] == 61524 && 
b[61525] == 61525 && 
b[61526] == 61526 && 
b[61527] == 61527 && 
b[61528] == 61528 && 
b[61529] == 61529 && 
b[61530] == 61530 && 
b[61531] == 61531 && 
b[61532] == 61532 && 
b[61533] == 61533 && 
b[61534] == 61534 && 
b[61535] == 61535 && 
b[61536] == 61536 && 
b[61537] == 61537 && 
b[61538] == 61538 && 
b[61539] == 61539 && 
b[61540] == 61540 && 
b[61541] == 61541 && 
b[61542] == 61542 && 
b[61543] == 61543 && 
b[61544] == 61544 && 
b[61545] == 61545 && 
b[61546] == 61546 && 
b[61547] == 61547 && 
b[61548] == 61548 && 
b[61549] == 61549 && 
b[61550] == 61550 && 
b[61551] == 61551 && 
b[61552] == 61552 && 
b[61553] == 61553 && 
b[61554] == 61554 && 
b[61555] == 61555 && 
b[61556] == 61556 && 
b[61557] == 61557 && 
b[61558] == 61558 && 
b[61559] == 61559 && 
b[61560] == 61560 && 
b[61561] == 61561 && 
b[61562] == 61562 && 
b[61563] == 61563 && 
b[61564] == 61564 && 
b[61565] == 61565 && 
b[61566] == 61566 && 
b[61567] == 61567 && 
b[61568] == 61568 && 
b[61569] == 61569 && 
b[61570] == 61570 && 
b[61571] == 61571 && 
b[61572] == 61572 && 
b[61573] == 61573 && 
b[61574] == 61574 && 
b[61575] == 61575 && 
b[61576] == 61576 && 
b[61577] == 61577 && 
b[61578] == 61578 && 
b[61579] == 61579 && 
b[61580] == 61580 && 
b[61581] == 61581 && 
b[61582] == 61582 && 
b[61583] == 61583 && 
b[61584] == 61584 && 
b[61585] == 61585 && 
b[61586] == 61586 && 
b[61587] == 61587 && 
b[61588] == 61588 && 
b[61589] == 61589 && 
b[61590] == 61590 && 
b[61591] == 61591 && 
b[61592] == 61592 && 
b[61593] == 61593 && 
b[61594] == 61594 && 
b[61595] == 61595 && 
b[61596] == 61596 && 
b[61597] == 61597 && 
b[61598] == 61598 && 
b[61599] == 61599 && 
b[61600] == 61600 && 
b[61601] == 61601 && 
b[61602] == 61602 && 
b[61603] == 61603 && 
b[61604] == 61604 && 
b[61605] == 61605 && 
b[61606] == 61606 && 
b[61607] == 61607 && 
b[61608] == 61608 && 
b[61609] == 61609 && 
b[61610] == 61610 && 
b[61611] == 61611 && 
b[61612] == 61612 && 
b[61613] == 61613 && 
b[61614] == 61614 && 
b[61615] == 61615 && 
b[61616] == 61616 && 
b[61617] == 61617 && 
b[61618] == 61618 && 
b[61619] == 61619 && 
b[61620] == 61620 && 
b[61621] == 61621 && 
b[61622] == 61622 && 
b[61623] == 61623 && 
b[61624] == 61624 && 
b[61625] == 61625 && 
b[61626] == 61626 && 
b[61627] == 61627 && 
b[61628] == 61628 && 
b[61629] == 61629 && 
b[61630] == 61630 && 
b[61631] == 61631 && 
b[61632] == 61632 && 
b[61633] == 61633 && 
b[61634] == 61634 && 
b[61635] == 61635 && 
b[61636] == 61636 && 
b[61637] == 61637 && 
b[61638] == 61638 && 
b[61639] == 61639 && 
b[61640] == 61640 && 
b[61641] == 61641 && 
b[61642] == 61642 && 
b[61643] == 61643 && 
b[61644] == 61644 && 
b[61645] == 61645 && 
b[61646] == 61646 && 
b[61647] == 61647 && 
b[61648] == 61648 && 
b[61649] == 61649 && 
b[61650] == 61650 && 
b[61651] == 61651 && 
b[61652] == 61652 && 
b[61653] == 61653 && 
b[61654] == 61654 && 
b[61655] == 61655 && 
b[61656] == 61656 && 
b[61657] == 61657 && 
b[61658] == 61658 && 
b[61659] == 61659 && 
b[61660] == 61660 && 
b[61661] == 61661 && 
b[61662] == 61662 && 
b[61663] == 61663 && 
b[61664] == 61664 && 
b[61665] == 61665 && 
b[61666] == 61666 && 
b[61667] == 61667 && 
b[61668] == 61668 && 
b[61669] == 61669 && 
b[61670] == 61670 && 
b[61671] == 61671 && 
b[61672] == 61672 && 
b[61673] == 61673 && 
b[61674] == 61674 && 
b[61675] == 61675 && 
b[61676] == 61676 && 
b[61677] == 61677 && 
b[61678] == 61678 && 
b[61679] == 61679 && 
b[61680] == 61680 && 
b[61681] == 61681 && 
b[61682] == 61682 && 
b[61683] == 61683 && 
b[61684] == 61684 && 
b[61685] == 61685 && 
b[61686] == 61686 && 
b[61687] == 61687 && 
b[61688] == 61688 && 
b[61689] == 61689 && 
b[61690] == 61690 && 
b[61691] == 61691 && 
b[61692] == 61692 && 
b[61693] == 61693 && 
b[61694] == 61694 && 
b[61695] == 61695 && 
b[61696] == 61696 && 
b[61697] == 61697 && 
b[61698] == 61698 && 
b[61699] == 61699 && 
b[61700] == 61700 && 
b[61701] == 61701 && 
b[61702] == 61702 && 
b[61703] == 61703 && 
b[61704] == 61704 && 
b[61705] == 61705 && 
b[61706] == 61706 && 
b[61707] == 61707 && 
b[61708] == 61708 && 
b[61709] == 61709 && 
b[61710] == 61710 && 
b[61711] == 61711 && 
b[61712] == 61712 && 
b[61713] == 61713 && 
b[61714] == 61714 && 
b[61715] == 61715 && 
b[61716] == 61716 && 
b[61717] == 61717 && 
b[61718] == 61718 && 
b[61719] == 61719 && 
b[61720] == 61720 && 
b[61721] == 61721 && 
b[61722] == 61722 && 
b[61723] == 61723 && 
b[61724] == 61724 && 
b[61725] == 61725 && 
b[61726] == 61726 && 
b[61727] == 61727 && 
b[61728] == 61728 && 
b[61729] == 61729 && 
b[61730] == 61730 && 
b[61731] == 61731 && 
b[61732] == 61732 && 
b[61733] == 61733 && 
b[61734] == 61734 && 
b[61735] == 61735 && 
b[61736] == 61736 && 
b[61737] == 61737 && 
b[61738] == 61738 && 
b[61739] == 61739 && 
b[61740] == 61740 && 
b[61741] == 61741 && 
b[61742] == 61742 && 
b[61743] == 61743 && 
b[61744] == 61744 && 
b[61745] == 61745 && 
b[61746] == 61746 && 
b[61747] == 61747 && 
b[61748] == 61748 && 
b[61749] == 61749 && 
b[61750] == 61750 && 
b[61751] == 61751 && 
b[61752] == 61752 && 
b[61753] == 61753 && 
b[61754] == 61754 && 
b[61755] == 61755 && 
b[61756] == 61756 && 
b[61757] == 61757 && 
b[61758] == 61758 && 
b[61759] == 61759 && 
b[61760] == 61760 && 
b[61761] == 61761 && 
b[61762] == 61762 && 
b[61763] == 61763 && 
b[61764] == 61764 && 
b[61765] == 61765 && 
b[61766] == 61766 && 
b[61767] == 61767 && 
b[61768] == 61768 && 
b[61769] == 61769 && 
b[61770] == 61770 && 
b[61771] == 61771 && 
b[61772] == 61772 && 
b[61773] == 61773 && 
b[61774] == 61774 && 
b[61775] == 61775 && 
b[61776] == 61776 && 
b[61777] == 61777 && 
b[61778] == 61778 && 
b[61779] == 61779 && 
b[61780] == 61780 && 
b[61781] == 61781 && 
b[61782] == 61782 && 
b[61783] == 61783 && 
b[61784] == 61784 && 
b[61785] == 61785 && 
b[61786] == 61786 && 
b[61787] == 61787 && 
b[61788] == 61788 && 
b[61789] == 61789 && 
b[61790] == 61790 && 
b[61791] == 61791 && 
b[61792] == 61792 && 
b[61793] == 61793 && 
b[61794] == 61794 && 
b[61795] == 61795 && 
b[61796] == 61796 && 
b[61797] == 61797 && 
b[61798] == 61798 && 
b[61799] == 61799 && 
b[61800] == 61800 && 
b[61801] == 61801 && 
b[61802] == 61802 && 
b[61803] == 61803 && 
b[61804] == 61804 && 
b[61805] == 61805 && 
b[61806] == 61806 && 
b[61807] == 61807 && 
b[61808] == 61808 && 
b[61809] == 61809 && 
b[61810] == 61810 && 
b[61811] == 61811 && 
b[61812] == 61812 && 
b[61813] == 61813 && 
b[61814] == 61814 && 
b[61815] == 61815 && 
b[61816] == 61816 && 
b[61817] == 61817 && 
b[61818] == 61818 && 
b[61819] == 61819 && 
b[61820] == 61820 && 
b[61821] == 61821 && 
b[61822] == 61822 && 
b[61823] == 61823 && 
b[61824] == 61824 && 
b[61825] == 61825 && 
b[61826] == 61826 && 
b[61827] == 61827 && 
b[61828] == 61828 && 
b[61829] == 61829 && 
b[61830] == 61830 && 
b[61831] == 61831 && 
b[61832] == 61832 && 
b[61833] == 61833 && 
b[61834] == 61834 && 
b[61835] == 61835 && 
b[61836] == 61836 && 
b[61837] == 61837 && 
b[61838] == 61838 && 
b[61839] == 61839 && 
b[61840] == 61840 && 
b[61841] == 61841 && 
b[61842] == 61842 && 
b[61843] == 61843 && 
b[61844] == 61844 && 
b[61845] == 61845 && 
b[61846] == 61846 && 
b[61847] == 61847 && 
b[61848] == 61848 && 
b[61849] == 61849 && 
b[61850] == 61850 && 
b[61851] == 61851 && 
b[61852] == 61852 && 
b[61853] == 61853 && 
b[61854] == 61854 && 
b[61855] == 61855 && 
b[61856] == 61856 && 
b[61857] == 61857 && 
b[61858] == 61858 && 
b[61859] == 61859 && 
b[61860] == 61860 && 
b[61861] == 61861 && 
b[61862] == 61862 && 
b[61863] == 61863 && 
b[61864] == 61864 && 
b[61865] == 61865 && 
b[61866] == 61866 && 
b[61867] == 61867 && 
b[61868] == 61868 && 
b[61869] == 61869 && 
b[61870] == 61870 && 
b[61871] == 61871 && 
b[61872] == 61872 && 
b[61873] == 61873 && 
b[61874] == 61874 && 
b[61875] == 61875 && 
b[61876] == 61876 && 
b[61877] == 61877 && 
b[61878] == 61878 && 
b[61879] == 61879 && 
b[61880] == 61880 && 
b[61881] == 61881 && 
b[61882] == 61882 && 
b[61883] == 61883 && 
b[61884] == 61884 && 
b[61885] == 61885 && 
b[61886] == 61886 && 
b[61887] == 61887 && 
b[61888] == 61888 && 
b[61889] == 61889 && 
b[61890] == 61890 && 
b[61891] == 61891 && 
b[61892] == 61892 && 
b[61893] == 61893 && 
b[61894] == 61894 && 
b[61895] == 61895 && 
b[61896] == 61896 && 
b[61897] == 61897 && 
b[61898] == 61898 && 
b[61899] == 61899 && 
b[61900] == 61900 && 
b[61901] == 61901 && 
b[61902] == 61902 && 
b[61903] == 61903 && 
b[61904] == 61904 && 
b[61905] == 61905 && 
b[61906] == 61906 && 
b[61907] == 61907 && 
b[61908] == 61908 && 
b[61909] == 61909 && 
b[61910] == 61910 && 
b[61911] == 61911 && 
b[61912] == 61912 && 
b[61913] == 61913 && 
b[61914] == 61914 && 
b[61915] == 61915 && 
b[61916] == 61916 && 
b[61917] == 61917 && 
b[61918] == 61918 && 
b[61919] == 61919 && 
b[61920] == 61920 && 
b[61921] == 61921 && 
b[61922] == 61922 && 
b[61923] == 61923 && 
b[61924] == 61924 && 
b[61925] == 61925 && 
b[61926] == 61926 && 
b[61927] == 61927 && 
b[61928] == 61928 && 
b[61929] == 61929 && 
b[61930] == 61930 && 
b[61931] == 61931 && 
b[61932] == 61932 && 
b[61933] == 61933 && 
b[61934] == 61934 && 
b[61935] == 61935 && 
b[61936] == 61936 && 
b[61937] == 61937 && 
b[61938] == 61938 && 
b[61939] == 61939 && 
b[61940] == 61940 && 
b[61941] == 61941 && 
b[61942] == 61942 && 
b[61943] == 61943 && 
b[61944] == 61944 && 
b[61945] == 61945 && 
b[61946] == 61946 && 
b[61947] == 61947 && 
b[61948] == 61948 && 
b[61949] == 61949 && 
b[61950] == 61950 && 
b[61951] == 61951 && 
b[61952] == 61952 && 
b[61953] == 61953 && 
b[61954] == 61954 && 
b[61955] == 61955 && 
b[61956] == 61956 && 
b[61957] == 61957 && 
b[61958] == 61958 && 
b[61959] == 61959 && 
b[61960] == 61960 && 
b[61961] == 61961 && 
b[61962] == 61962 && 
b[61963] == 61963 && 
b[61964] == 61964 && 
b[61965] == 61965 && 
b[61966] == 61966 && 
b[61967] == 61967 && 
b[61968] == 61968 && 
b[61969] == 61969 && 
b[61970] == 61970 && 
b[61971] == 61971 && 
b[61972] == 61972 && 
b[61973] == 61973 && 
b[61974] == 61974 && 
b[61975] == 61975 && 
b[61976] == 61976 && 
b[61977] == 61977 && 
b[61978] == 61978 && 
b[61979] == 61979 && 
b[61980] == 61980 && 
b[61981] == 61981 && 
b[61982] == 61982 && 
b[61983] == 61983 && 
b[61984] == 61984 && 
b[61985] == 61985 && 
b[61986] == 61986 && 
b[61987] == 61987 && 
b[61988] == 61988 && 
b[61989] == 61989 && 
b[61990] == 61990 && 
b[61991] == 61991 && 
b[61992] == 61992 && 
b[61993] == 61993 && 
b[61994] == 61994 && 
b[61995] == 61995 && 
b[61996] == 61996 && 
b[61997] == 61997 && 
b[61998] == 61998 && 
b[61999] == 61999 && 
b[62000] == 62000 && 
b[62001] == 62001 && 
b[62002] == 62002 && 
b[62003] == 62003 && 
b[62004] == 62004 && 
b[62005] == 62005 && 
b[62006] == 62006 && 
b[62007] == 62007 && 
b[62008] == 62008 && 
b[62009] == 62009 && 
b[62010] == 62010 && 
b[62011] == 62011 && 
b[62012] == 62012 && 
b[62013] == 62013 && 
b[62014] == 62014 && 
b[62015] == 62015 && 
b[62016] == 62016 && 
b[62017] == 62017 && 
b[62018] == 62018 && 
b[62019] == 62019 && 
b[62020] == 62020 && 
b[62021] == 62021 && 
b[62022] == 62022 && 
b[62023] == 62023 && 
b[62024] == 62024 && 
b[62025] == 62025 && 
b[62026] == 62026 && 
b[62027] == 62027 && 
b[62028] == 62028 && 
b[62029] == 62029 && 
b[62030] == 62030 && 
b[62031] == 62031 && 
b[62032] == 62032 && 
b[62033] == 62033 && 
b[62034] == 62034 && 
b[62035] == 62035 && 
b[62036] == 62036 && 
b[62037] == 62037 && 
b[62038] == 62038 && 
b[62039] == 62039 && 
b[62040] == 62040 && 
b[62041] == 62041 && 
b[62042] == 62042 && 
b[62043] == 62043 && 
b[62044] == 62044 && 
b[62045] == 62045 && 
b[62046] == 62046 && 
b[62047] == 62047 && 
b[62048] == 62048 && 
b[62049] == 62049 && 
b[62050] == 62050 && 
b[62051] == 62051 && 
b[62052] == 62052 && 
b[62053] == 62053 && 
b[62054] == 62054 && 
b[62055] == 62055 && 
b[62056] == 62056 && 
b[62057] == 62057 && 
b[62058] == 62058 && 
b[62059] == 62059 && 
b[62060] == 62060 && 
b[62061] == 62061 && 
b[62062] == 62062 && 
b[62063] == 62063 && 
b[62064] == 62064 && 
b[62065] == 62065 && 
b[62066] == 62066 && 
b[62067] == 62067 && 
b[62068] == 62068 && 
b[62069] == 62069 && 
b[62070] == 62070 && 
b[62071] == 62071 && 
b[62072] == 62072 && 
b[62073] == 62073 && 
b[62074] == 62074 && 
b[62075] == 62075 && 
b[62076] == 62076 && 
b[62077] == 62077 && 
b[62078] == 62078 && 
b[62079] == 62079 && 
b[62080] == 62080 && 
b[62081] == 62081 && 
b[62082] == 62082 && 
b[62083] == 62083 && 
b[62084] == 62084 && 
b[62085] == 62085 && 
b[62086] == 62086 && 
b[62087] == 62087 && 
b[62088] == 62088 && 
b[62089] == 62089 && 
b[62090] == 62090 && 
b[62091] == 62091 && 
b[62092] == 62092 && 
b[62093] == 62093 && 
b[62094] == 62094 && 
b[62095] == 62095 && 
b[62096] == 62096 && 
b[62097] == 62097 && 
b[62098] == 62098 && 
b[62099] == 62099 && 
b[62100] == 62100 && 
b[62101] == 62101 && 
b[62102] == 62102 && 
b[62103] == 62103 && 
b[62104] == 62104 && 
b[62105] == 62105 && 
b[62106] == 62106 && 
b[62107] == 62107 && 
b[62108] == 62108 && 
b[62109] == 62109 && 
b[62110] == 62110 && 
b[62111] == 62111 && 
b[62112] == 62112 && 
b[62113] == 62113 && 
b[62114] == 62114 && 
b[62115] == 62115 && 
b[62116] == 62116 && 
b[62117] == 62117 && 
b[62118] == 62118 && 
b[62119] == 62119 && 
b[62120] == 62120 && 
b[62121] == 62121 && 
b[62122] == 62122 && 
b[62123] == 62123 && 
b[62124] == 62124 && 
b[62125] == 62125 && 
b[62126] == 62126 && 
b[62127] == 62127 && 
b[62128] == 62128 && 
b[62129] == 62129 && 
b[62130] == 62130 && 
b[62131] == 62131 && 
b[62132] == 62132 && 
b[62133] == 62133 && 
b[62134] == 62134 && 
b[62135] == 62135 && 
b[62136] == 62136 && 
b[62137] == 62137 && 
b[62138] == 62138 && 
b[62139] == 62139 && 
b[62140] == 62140 && 
b[62141] == 62141 && 
b[62142] == 62142 && 
b[62143] == 62143 && 
b[62144] == 62144 && 
b[62145] == 62145 && 
b[62146] == 62146 && 
b[62147] == 62147 && 
b[62148] == 62148 && 
b[62149] == 62149 && 
b[62150] == 62150 && 
b[62151] == 62151 && 
b[62152] == 62152 && 
b[62153] == 62153 && 
b[62154] == 62154 && 
b[62155] == 62155 && 
b[62156] == 62156 && 
b[62157] == 62157 && 
b[62158] == 62158 && 
b[62159] == 62159 && 
b[62160] == 62160 && 
b[62161] == 62161 && 
b[62162] == 62162 && 
b[62163] == 62163 && 
b[62164] == 62164 && 
b[62165] == 62165 && 
b[62166] == 62166 && 
b[62167] == 62167 && 
b[62168] == 62168 && 
b[62169] == 62169 && 
b[62170] == 62170 && 
b[62171] == 62171 && 
b[62172] == 62172 && 
b[62173] == 62173 && 
b[62174] == 62174 && 
b[62175] == 62175 && 
b[62176] == 62176 && 
b[62177] == 62177 && 
b[62178] == 62178 && 
b[62179] == 62179 && 
b[62180] == 62180 && 
b[62181] == 62181 && 
b[62182] == 62182 && 
b[62183] == 62183 && 
b[62184] == 62184 && 
b[62185] == 62185 && 
b[62186] == 62186 && 
b[62187] == 62187 && 
b[62188] == 62188 && 
b[62189] == 62189 && 
b[62190] == 62190 && 
b[62191] == 62191 && 
b[62192] == 62192 && 
b[62193] == 62193 && 
b[62194] == 62194 && 
b[62195] == 62195 && 
b[62196] == 62196 && 
b[62197] == 62197 && 
b[62198] == 62198 && 
b[62199] == 62199 && 
b[62200] == 62200 && 
b[62201] == 62201 && 
b[62202] == 62202 && 
b[62203] == 62203 && 
b[62204] == 62204 && 
b[62205] == 62205 && 
b[62206] == 62206 && 
b[62207] == 62207 && 
b[62208] == 62208 && 
b[62209] == 62209 && 
b[62210] == 62210 && 
b[62211] == 62211 && 
b[62212] == 62212 && 
b[62213] == 62213 && 
b[62214] == 62214 && 
b[62215] == 62215 && 
b[62216] == 62216 && 
b[62217] == 62217 && 
b[62218] == 62218 && 
b[62219] == 62219 && 
b[62220] == 62220 && 
b[62221] == 62221 && 
b[62222] == 62222 && 
b[62223] == 62223 && 
b[62224] == 62224 && 
b[62225] == 62225 && 
b[62226] == 62226 && 
b[62227] == 62227 && 
b[62228] == 62228 && 
b[62229] == 62229 && 
b[62230] == 62230 && 
b[62231] == 62231 && 
b[62232] == 62232 && 
b[62233] == 62233 && 
b[62234] == 62234 && 
b[62235] == 62235 && 
b[62236] == 62236 && 
b[62237] == 62237 && 
b[62238] == 62238 && 
b[62239] == 62239 && 
b[62240] == 62240 && 
b[62241] == 62241 && 
b[62242] == 62242 && 
b[62243] == 62243 && 
b[62244] == 62244 && 
b[62245] == 62245 && 
b[62246] == 62246 && 
b[62247] == 62247 && 
b[62248] == 62248 && 
b[62249] == 62249 && 
b[62250] == 62250 && 
b[62251] == 62251 && 
b[62252] == 62252 && 
b[62253] == 62253 && 
b[62254] == 62254 && 
b[62255] == 62255 && 
b[62256] == 62256 && 
b[62257] == 62257 && 
b[62258] == 62258 && 
b[62259] == 62259 && 
b[62260] == 62260 && 
b[62261] == 62261 && 
b[62262] == 62262 && 
b[62263] == 62263 && 
b[62264] == 62264 && 
b[62265] == 62265 && 
b[62266] == 62266 && 
b[62267] == 62267 && 
b[62268] == 62268 && 
b[62269] == 62269 && 
b[62270] == 62270 && 
b[62271] == 62271 && 
b[62272] == 62272 && 
b[62273] == 62273 && 
b[62274] == 62274 && 
b[62275] == 62275 && 
b[62276] == 62276 && 
b[62277] == 62277 && 
b[62278] == 62278 && 
b[62279] == 62279 && 
b[62280] == 62280 && 
b[62281] == 62281 && 
b[62282] == 62282 && 
b[62283] == 62283 && 
b[62284] == 62284 && 
b[62285] == 62285 && 
b[62286] == 62286 && 
b[62287] == 62287 && 
b[62288] == 62288 && 
b[62289] == 62289 && 
b[62290] == 62290 && 
b[62291] == 62291 && 
b[62292] == 62292 && 
b[62293] == 62293 && 
b[62294] == 62294 && 
b[62295] == 62295 && 
b[62296] == 62296 && 
b[62297] == 62297 && 
b[62298] == 62298 && 
b[62299] == 62299 && 
b[62300] == 62300 && 
b[62301] == 62301 && 
b[62302] == 62302 && 
b[62303] == 62303 && 
b[62304] == 62304 && 
b[62305] == 62305 && 
b[62306] == 62306 && 
b[62307] == 62307 && 
b[62308] == 62308 && 
b[62309] == 62309 && 
b[62310] == 62310 && 
b[62311] == 62311 && 
b[62312] == 62312 && 
b[62313] == 62313 && 
b[62314] == 62314 && 
b[62315] == 62315 && 
b[62316] == 62316 && 
b[62317] == 62317 && 
b[62318] == 62318 && 
b[62319] == 62319 && 
b[62320] == 62320 && 
b[62321] == 62321 && 
b[62322] == 62322 && 
b[62323] == 62323 && 
b[62324] == 62324 && 
b[62325] == 62325 && 
b[62326] == 62326 && 
b[62327] == 62327 && 
b[62328] == 62328 && 
b[62329] == 62329 && 
b[62330] == 62330 && 
b[62331] == 62331 && 
b[62332] == 62332 && 
b[62333] == 62333 && 
b[62334] == 62334 && 
b[62335] == 62335 && 
b[62336] == 62336 && 
b[62337] == 62337 && 
b[62338] == 62338 && 
b[62339] == 62339 && 
b[62340] == 62340 && 
b[62341] == 62341 && 
b[62342] == 62342 && 
b[62343] == 62343 && 
b[62344] == 62344 && 
b[62345] == 62345 && 
b[62346] == 62346 && 
b[62347] == 62347 && 
b[62348] == 62348 && 
b[62349] == 62349 && 
b[62350] == 62350 && 
b[62351] == 62351 && 
b[62352] == 62352 && 
b[62353] == 62353 && 
b[62354] == 62354 && 
b[62355] == 62355 && 
b[62356] == 62356 && 
b[62357] == 62357 && 
b[62358] == 62358 && 
b[62359] == 62359 && 
b[62360] == 62360 && 
b[62361] == 62361 && 
b[62362] == 62362 && 
b[62363] == 62363 && 
b[62364] == 62364 && 
b[62365] == 62365 && 
b[62366] == 62366 && 
b[62367] == 62367 && 
b[62368] == 62368 && 
b[62369] == 62369 && 
b[62370] == 62370 && 
b[62371] == 62371 && 
b[62372] == 62372 && 
b[62373] == 62373 && 
b[62374] == 62374 && 
b[62375] == 62375 && 
b[62376] == 62376 && 
b[62377] == 62377 && 
b[62378] == 62378 && 
b[62379] == 62379 && 
b[62380] == 62380 && 
b[62381] == 62381 && 
b[62382] == 62382 && 
b[62383] == 62383 && 
b[62384] == 62384 && 
b[62385] == 62385 && 
b[62386] == 62386 && 
b[62387] == 62387 && 
b[62388] == 62388 && 
b[62389] == 62389 && 
b[62390] == 62390 && 
b[62391] == 62391 && 
b[62392] == 62392 && 
b[62393] == 62393 && 
b[62394] == 62394 && 
b[62395] == 62395 && 
b[62396] == 62396 && 
b[62397] == 62397 && 
b[62398] == 62398 && 
b[62399] == 62399 && 
b[62400] == 62400 && 
b[62401] == 62401 && 
b[62402] == 62402 && 
b[62403] == 62403 && 
b[62404] == 62404 && 
b[62405] == 62405 && 
b[62406] == 62406 && 
b[62407] == 62407 && 
b[62408] == 62408 && 
b[62409] == 62409 && 
b[62410] == 62410 && 
b[62411] == 62411 && 
b[62412] == 62412 && 
b[62413] == 62413 && 
b[62414] == 62414 && 
b[62415] == 62415 && 
b[62416] == 62416 && 
b[62417] == 62417 && 
b[62418] == 62418 && 
b[62419] == 62419 && 
b[62420] == 62420 && 
b[62421] == 62421 && 
b[62422] == 62422 && 
b[62423] == 62423 && 
b[62424] == 62424 && 
b[62425] == 62425 && 
b[62426] == 62426 && 
b[62427] == 62427 && 
b[62428] == 62428 && 
b[62429] == 62429 && 
b[62430] == 62430 && 
b[62431] == 62431 && 
b[62432] == 62432 && 
b[62433] == 62433 && 
b[62434] == 62434 && 
b[62435] == 62435 && 
b[62436] == 62436 && 
b[62437] == 62437 && 
b[62438] == 62438 && 
b[62439] == 62439 && 
b[62440] == 62440 && 
b[62441] == 62441 && 
b[62442] == 62442 && 
b[62443] == 62443 && 
b[62444] == 62444 && 
b[62445] == 62445 && 
b[62446] == 62446 && 
b[62447] == 62447 && 
b[62448] == 62448 && 
b[62449] == 62449 && 
b[62450] == 62450 && 
b[62451] == 62451 && 
b[62452] == 62452 && 
b[62453] == 62453 && 
b[62454] == 62454 && 
b[62455] == 62455 && 
b[62456] == 62456 && 
b[62457] == 62457 && 
b[62458] == 62458 && 
b[62459] == 62459 && 
b[62460] == 62460 && 
b[62461] == 62461 && 
b[62462] == 62462 && 
b[62463] == 62463 && 
b[62464] == 62464 && 
b[62465] == 62465 && 
b[62466] == 62466 && 
b[62467] == 62467 && 
b[62468] == 62468 && 
b[62469] == 62469 && 
b[62470] == 62470 && 
b[62471] == 62471 && 
b[62472] == 62472 && 
b[62473] == 62473 && 
b[62474] == 62474 && 
b[62475] == 62475 && 
b[62476] == 62476 && 
b[62477] == 62477 && 
b[62478] == 62478 && 
b[62479] == 62479 && 
b[62480] == 62480 && 
b[62481] == 62481 && 
b[62482] == 62482 && 
b[62483] == 62483 && 
b[62484] == 62484 && 
b[62485] == 62485 && 
b[62486] == 62486 && 
b[62487] == 62487 && 
b[62488] == 62488 && 
b[62489] == 62489 && 
b[62490] == 62490 && 
b[62491] == 62491 && 
b[62492] == 62492 && 
b[62493] == 62493 && 
b[62494] == 62494 && 
b[62495] == 62495 && 
b[62496] == 62496 && 
b[62497] == 62497 && 
b[62498] == 62498 && 
b[62499] == 62499 && 
b[62500] == 62500 && 
b[62501] == 62501 && 
b[62502] == 62502 && 
b[62503] == 62503 && 
b[62504] == 62504 && 
b[62505] == 62505 && 
b[62506] == 62506 && 
b[62507] == 62507 && 
b[62508] == 62508 && 
b[62509] == 62509 && 
b[62510] == 62510 && 
b[62511] == 62511 && 
b[62512] == 62512 && 
b[62513] == 62513 && 
b[62514] == 62514 && 
b[62515] == 62515 && 
b[62516] == 62516 && 
b[62517] == 62517 && 
b[62518] == 62518 && 
b[62519] == 62519 && 
b[62520] == 62520 && 
b[62521] == 62521 && 
b[62522] == 62522 && 
b[62523] == 62523 && 
b[62524] == 62524 && 
b[62525] == 62525 && 
b[62526] == 62526 && 
b[62527] == 62527 && 
b[62528] == 62528 && 
b[62529] == 62529 && 
b[62530] == 62530 && 
b[62531] == 62531 && 
b[62532] == 62532 && 
b[62533] == 62533 && 
b[62534] == 62534 && 
b[62535] == 62535 && 
b[62536] == 62536 && 
b[62537] == 62537 && 
b[62538] == 62538 && 
b[62539] == 62539 && 
b[62540] == 62540 && 
b[62541] == 62541 && 
b[62542] == 62542 && 
b[62543] == 62543 && 
b[62544] == 62544 && 
b[62545] == 62545 && 
b[62546] == 62546 && 
b[62547] == 62547 && 
b[62548] == 62548 && 
b[62549] == 62549 && 
b[62550] == 62550 && 
b[62551] == 62551 && 
b[62552] == 62552 && 
b[62553] == 62553 && 
b[62554] == 62554 && 
b[62555] == 62555 && 
b[62556] == 62556 && 
b[62557] == 62557 && 
b[62558] == 62558 && 
b[62559] == 62559 && 
b[62560] == 62560 && 
b[62561] == 62561 && 
b[62562] == 62562 && 
b[62563] == 62563 && 
b[62564] == 62564 && 
b[62565] == 62565 && 
b[62566] == 62566 && 
b[62567] == 62567 && 
b[62568] == 62568 && 
b[62569] == 62569 && 
b[62570] == 62570 && 
b[62571] == 62571 && 
b[62572] == 62572 && 
b[62573] == 62573 && 
b[62574] == 62574 && 
b[62575] == 62575 && 
b[62576] == 62576 && 
b[62577] == 62577 && 
b[62578] == 62578 && 
b[62579] == 62579 && 
b[62580] == 62580 && 
b[62581] == 62581 && 
b[62582] == 62582 && 
b[62583] == 62583 && 
b[62584] == 62584 && 
b[62585] == 62585 && 
b[62586] == 62586 && 
b[62587] == 62587 && 
b[62588] == 62588 && 
b[62589] == 62589 && 
b[62590] == 62590 && 
b[62591] == 62591 && 
b[62592] == 62592 && 
b[62593] == 62593 && 
b[62594] == 62594 && 
b[62595] == 62595 && 
b[62596] == 62596 && 
b[62597] == 62597 && 
b[62598] == 62598 && 
b[62599] == 62599 && 
b[62600] == 62600 && 
b[62601] == 62601 && 
b[62602] == 62602 && 
b[62603] == 62603 && 
b[62604] == 62604 && 
b[62605] == 62605 && 
b[62606] == 62606 && 
b[62607] == 62607 && 
b[62608] == 62608 && 
b[62609] == 62609 && 
b[62610] == 62610 && 
b[62611] == 62611 && 
b[62612] == 62612 && 
b[62613] == 62613 && 
b[62614] == 62614 && 
b[62615] == 62615 && 
b[62616] == 62616 && 
b[62617] == 62617 && 
b[62618] == 62618 && 
b[62619] == 62619 && 
b[62620] == 62620 && 
b[62621] == 62621 && 
b[62622] == 62622 && 
b[62623] == 62623 && 
b[62624] == 62624 && 
b[62625] == 62625 && 
b[62626] == 62626 && 
b[62627] == 62627 && 
b[62628] == 62628 && 
b[62629] == 62629 && 
b[62630] == 62630 && 
b[62631] == 62631 && 
b[62632] == 62632 && 
b[62633] == 62633 && 
b[62634] == 62634 && 
b[62635] == 62635 && 
b[62636] == 62636 && 
b[62637] == 62637 && 
b[62638] == 62638 && 
b[62639] == 62639 && 
b[62640] == 62640 && 
b[62641] == 62641 && 
b[62642] == 62642 && 
b[62643] == 62643 && 
b[62644] == 62644 && 
b[62645] == 62645 && 
b[62646] == 62646 && 
b[62647] == 62647 && 
b[62648] == 62648 && 
b[62649] == 62649 && 
b[62650] == 62650 && 
b[62651] == 62651 && 
b[62652] == 62652 && 
b[62653] == 62653 && 
b[62654] == 62654 && 
b[62655] == 62655 && 
b[62656] == 62656 && 
b[62657] == 62657 && 
b[62658] == 62658 && 
b[62659] == 62659 && 
b[62660] == 62660 && 
b[62661] == 62661 && 
b[62662] == 62662 && 
b[62663] == 62663 && 
b[62664] == 62664 && 
b[62665] == 62665 && 
b[62666] == 62666 && 
b[62667] == 62667 && 
b[62668] == 62668 && 
b[62669] == 62669 && 
b[62670] == 62670 && 
b[62671] == 62671 && 
b[62672] == 62672 && 
b[62673] == 62673 && 
b[62674] == 62674 && 
b[62675] == 62675 && 
b[62676] == 62676 && 
b[62677] == 62677 && 
b[62678] == 62678 && 
b[62679] == 62679 && 
b[62680] == 62680 && 
b[62681] == 62681 && 
b[62682] == 62682 && 
b[62683] == 62683 && 
b[62684] == 62684 && 
b[62685] == 62685 && 
b[62686] == 62686 && 
b[62687] == 62687 && 
b[62688] == 62688 && 
b[62689] == 62689 && 
b[62690] == 62690 && 
b[62691] == 62691 && 
b[62692] == 62692 && 
b[62693] == 62693 && 
b[62694] == 62694 && 
b[62695] == 62695 && 
b[62696] == 62696 && 
b[62697] == 62697 && 
b[62698] == 62698 && 
b[62699] == 62699 && 
b[62700] == 62700 && 
b[62701] == 62701 && 
b[62702] == 62702 && 
b[62703] == 62703 && 
b[62704] == 62704 && 
b[62705] == 62705 && 
b[62706] == 62706 && 
b[62707] == 62707 && 
b[62708] == 62708 && 
b[62709] == 62709 && 
b[62710] == 62710 && 
b[62711] == 62711 && 
b[62712] == 62712 && 
b[62713] == 62713 && 
b[62714] == 62714 && 
b[62715] == 62715 && 
b[62716] == 62716 && 
b[62717] == 62717 && 
b[62718] == 62718 && 
b[62719] == 62719 && 
b[62720] == 62720 && 
b[62721] == 62721 && 
b[62722] == 62722 && 
b[62723] == 62723 && 
b[62724] == 62724 && 
b[62725] == 62725 && 
b[62726] == 62726 && 
b[62727] == 62727 && 
b[62728] == 62728 && 
b[62729] == 62729 && 
b[62730] == 62730 && 
b[62731] == 62731 && 
b[62732] == 62732 && 
b[62733] == 62733 && 
b[62734] == 62734 && 
b[62735] == 62735 && 
b[62736] == 62736 && 
b[62737] == 62737 && 
b[62738] == 62738 && 
b[62739] == 62739 && 
b[62740] == 62740 && 
b[62741] == 62741 && 
b[62742] == 62742 && 
b[62743] == 62743 && 
b[62744] == 62744 && 
b[62745] == 62745 && 
b[62746] == 62746 && 
b[62747] == 62747 && 
b[62748] == 62748 && 
b[62749] == 62749 && 
b[62750] == 62750 && 
b[62751] == 62751 && 
b[62752] == 62752 && 
b[62753] == 62753 && 
b[62754] == 62754 && 
b[62755] == 62755 && 
b[62756] == 62756 && 
b[62757] == 62757 && 
b[62758] == 62758 && 
b[62759] == 62759 && 
b[62760] == 62760 && 
b[62761] == 62761 && 
b[62762] == 62762 && 
b[62763] == 62763 && 
b[62764] == 62764 && 
b[62765] == 62765 && 
b[62766] == 62766 && 
b[62767] == 62767 && 
b[62768] == 62768 && 
b[62769] == 62769 && 
b[62770] == 62770 && 
b[62771] == 62771 && 
b[62772] == 62772 && 
b[62773] == 62773 && 
b[62774] == 62774 && 
b[62775] == 62775 && 
b[62776] == 62776 && 
b[62777] == 62777 && 
b[62778] == 62778 && 
b[62779] == 62779 && 
b[62780] == 62780 && 
b[62781] == 62781 && 
b[62782] == 62782 && 
b[62783] == 62783 && 
b[62784] == 62784 && 
b[62785] == 62785 && 
b[62786] == 62786 && 
b[62787] == 62787 && 
b[62788] == 62788 && 
b[62789] == 62789 && 
b[62790] == 62790 && 
b[62791] == 62791 && 
b[62792] == 62792 && 
b[62793] == 62793 && 
b[62794] == 62794 && 
b[62795] == 62795 && 
b[62796] == 62796 && 
b[62797] == 62797 && 
b[62798] == 62798 && 
b[62799] == 62799 && 
b[62800] == 62800 && 
b[62801] == 62801 && 
b[62802] == 62802 && 
b[62803] == 62803 && 
b[62804] == 62804 && 
b[62805] == 62805 && 
b[62806] == 62806 && 
b[62807] == 62807 && 
b[62808] == 62808 && 
b[62809] == 62809 && 
b[62810] == 62810 && 
b[62811] == 62811 && 
b[62812] == 62812 && 
b[62813] == 62813 && 
b[62814] == 62814 && 
b[62815] == 62815 && 
b[62816] == 62816 && 
b[62817] == 62817 && 
b[62818] == 62818 && 
b[62819] == 62819 && 
b[62820] == 62820 && 
b[62821] == 62821 && 
b[62822] == 62822 && 
b[62823] == 62823 && 
b[62824] == 62824 && 
b[62825] == 62825 && 
b[62826] == 62826 && 
b[62827] == 62827 && 
b[62828] == 62828 && 
b[62829] == 62829 && 
b[62830] == 62830 && 
b[62831] == 62831 && 
b[62832] == 62832 && 
b[62833] == 62833 && 
b[62834] == 62834 && 
b[62835] == 62835 && 
b[62836] == 62836 && 
b[62837] == 62837 && 
b[62838] == 62838 && 
b[62839] == 62839 && 
b[62840] == 62840 && 
b[62841] == 62841 && 
b[62842] == 62842 && 
b[62843] == 62843 && 
b[62844] == 62844 && 
b[62845] == 62845 && 
b[62846] == 62846 && 
b[62847] == 62847 && 
b[62848] == 62848 && 
b[62849] == 62849 && 
b[62850] == 62850 && 
b[62851] == 62851 && 
b[62852] == 62852 && 
b[62853] == 62853 && 
b[62854] == 62854 && 
b[62855] == 62855 && 
b[62856] == 62856 && 
b[62857] == 62857 && 
b[62858] == 62858 && 
b[62859] == 62859 && 
b[62860] == 62860 && 
b[62861] == 62861 && 
b[62862] == 62862 && 
b[62863] == 62863 && 
b[62864] == 62864 && 
b[62865] == 62865 && 
b[62866] == 62866 && 
b[62867] == 62867 && 
b[62868] == 62868 && 
b[62869] == 62869 && 
b[62870] == 62870 && 
b[62871] == 62871 && 
b[62872] == 62872 && 
b[62873] == 62873 && 
b[62874] == 62874 && 
b[62875] == 62875 && 
b[62876] == 62876 && 
b[62877] == 62877 && 
b[62878] == 62878 && 
b[62879] == 62879 && 
b[62880] == 62880 && 
b[62881] == 62881 && 
b[62882] == 62882 && 
b[62883] == 62883 && 
b[62884] == 62884 && 
b[62885] == 62885 && 
b[62886] == 62886 && 
b[62887] == 62887 && 
b[62888] == 62888 && 
b[62889] == 62889 && 
b[62890] == 62890 && 
b[62891] == 62891 && 
b[62892] == 62892 && 
b[62893] == 62893 && 
b[62894] == 62894 && 
b[62895] == 62895 && 
b[62896] == 62896 && 
b[62897] == 62897 && 
b[62898] == 62898 && 
b[62899] == 62899 && 
b[62900] == 62900 && 
b[62901] == 62901 && 
b[62902] == 62902 && 
b[62903] == 62903 && 
b[62904] == 62904 && 
b[62905] == 62905 && 
b[62906] == 62906 && 
b[62907] == 62907 && 
b[62908] == 62908 && 
b[62909] == 62909 && 
b[62910] == 62910 && 
b[62911] == 62911 && 
b[62912] == 62912 && 
b[62913] == 62913 && 
b[62914] == 62914 && 
b[62915] == 62915 && 
b[62916] == 62916 && 
b[62917] == 62917 && 
b[62918] == 62918 && 
b[62919] == 62919 && 
b[62920] == 62920 && 
b[62921] == 62921 && 
b[62922] == 62922 && 
b[62923] == 62923 && 
b[62924] == 62924 && 
b[62925] == 62925 && 
b[62926] == 62926 && 
b[62927] == 62927 && 
b[62928] == 62928 && 
b[62929] == 62929 && 
b[62930] == 62930 && 
b[62931] == 62931 && 
b[62932] == 62932 && 
b[62933] == 62933 && 
b[62934] == 62934 && 
b[62935] == 62935 && 
b[62936] == 62936 && 
b[62937] == 62937 && 
b[62938] == 62938 && 
b[62939] == 62939 && 
b[62940] == 62940 && 
b[62941] == 62941 && 
b[62942] == 62942 && 
b[62943] == 62943 && 
b[62944] == 62944 && 
b[62945] == 62945 && 
b[62946] == 62946 && 
b[62947] == 62947 && 
b[62948] == 62948 && 
b[62949] == 62949 && 
b[62950] == 62950 && 
b[62951] == 62951 && 
b[62952] == 62952 && 
b[62953] == 62953 && 
b[62954] == 62954 && 
b[62955] == 62955 && 
b[62956] == 62956 && 
b[62957] == 62957 && 
b[62958] == 62958 && 
b[62959] == 62959 && 
b[62960] == 62960 && 
b[62961] == 62961 && 
b[62962] == 62962 && 
b[62963] == 62963 && 
b[62964] == 62964 && 
b[62965] == 62965 && 
b[62966] == 62966 && 
b[62967] == 62967 && 
b[62968] == 62968 && 
b[62969] == 62969 && 
b[62970] == 62970 && 
b[62971] == 62971 && 
b[62972] == 62972 && 
b[62973] == 62973 && 
b[62974] == 62974 && 
b[62975] == 62975 && 
b[62976] == 62976 && 
b[62977] == 62977 && 
b[62978] == 62978 && 
b[62979] == 62979 && 
b[62980] == 62980 && 
b[62981] == 62981 && 
b[62982] == 62982 && 
b[62983] == 62983 && 
b[62984] == 62984 && 
b[62985] == 62985 && 
b[62986] == 62986 && 
b[62987] == 62987 && 
b[62988] == 62988 && 
b[62989] == 62989 && 
b[62990] == 62990 && 
b[62991] == 62991 && 
b[62992] == 62992 && 
b[62993] == 62993 && 
b[62994] == 62994 && 
b[62995] == 62995 && 
b[62996] == 62996 && 
b[62997] == 62997 && 
b[62998] == 62998 && 
b[62999] == 62999 && 
b[63000] == 63000 && 
b[63001] == 63001 && 
b[63002] == 63002 && 
b[63003] == 63003 && 
b[63004] == 63004 && 
b[63005] == 63005 && 
b[63006] == 63006 && 
b[63007] == 63007 && 
b[63008] == 63008 && 
b[63009] == 63009 && 
b[63010] == 63010 && 
b[63011] == 63011 && 
b[63012] == 63012 && 
b[63013] == 63013 && 
b[63014] == 63014 && 
b[63015] == 63015 && 
b[63016] == 63016 && 
b[63017] == 63017 && 
b[63018] == 63018 && 
b[63019] == 63019 && 
b[63020] == 63020 && 
b[63021] == 63021 && 
b[63022] == 63022 && 
b[63023] == 63023 && 
b[63024] == 63024 && 
b[63025] == 63025 && 
b[63026] == 63026 && 
b[63027] == 63027 && 
b[63028] == 63028 && 
b[63029] == 63029 && 
b[63030] == 63030 && 
b[63031] == 63031 && 
b[63032] == 63032 && 
b[63033] == 63033 && 
b[63034] == 63034 && 
b[63035] == 63035 && 
b[63036] == 63036 && 
b[63037] == 63037 && 
b[63038] == 63038 && 
b[63039] == 63039 && 
b[63040] == 63040 && 
b[63041] == 63041 && 
b[63042] == 63042 && 
b[63043] == 63043 && 
b[63044] == 63044 && 
b[63045] == 63045 && 
b[63046] == 63046 && 
b[63047] == 63047 && 
b[63048] == 63048 && 
b[63049] == 63049 && 
b[63050] == 63050 && 
b[63051] == 63051 && 
b[63052] == 63052 && 
b[63053] == 63053 && 
b[63054] == 63054 && 
b[63055] == 63055 && 
b[63056] == 63056 && 
b[63057] == 63057 && 
b[63058] == 63058 && 
b[63059] == 63059 && 
b[63060] == 63060 && 
b[63061] == 63061 && 
b[63062] == 63062 && 
b[63063] == 63063 && 
b[63064] == 63064 && 
b[63065] == 63065 && 
b[63066] == 63066 && 
b[63067] == 63067 && 
b[63068] == 63068 && 
b[63069] == 63069 && 
b[63070] == 63070 && 
b[63071] == 63071 && 
b[63072] == 63072 && 
b[63073] == 63073 && 
b[63074] == 63074 && 
b[63075] == 63075 && 
b[63076] == 63076 && 
b[63077] == 63077 && 
b[63078] == 63078 && 
b[63079] == 63079 && 
b[63080] == 63080 && 
b[63081] == 63081 && 
b[63082] == 63082 && 
b[63083] == 63083 && 
b[63084] == 63084 && 
b[63085] == 63085 && 
b[63086] == 63086 && 
b[63087] == 63087 && 
b[63088] == 63088 && 
b[63089] == 63089 && 
b[63090] == 63090 && 
b[63091] == 63091 && 
b[63092] == 63092 && 
b[63093] == 63093 && 
b[63094] == 63094 && 
b[63095] == 63095 && 
b[63096] == 63096 && 
b[63097] == 63097 && 
b[63098] == 63098 && 
b[63099] == 63099 && 
b[63100] == 63100 && 
b[63101] == 63101 && 
b[63102] == 63102 && 
b[63103] == 63103 && 
b[63104] == 63104 && 
b[63105] == 63105 && 
b[63106] == 63106 && 
b[63107] == 63107 && 
b[63108] == 63108 && 
b[63109] == 63109 && 
b[63110] == 63110 && 
b[63111] == 63111 && 
b[63112] == 63112 && 
b[63113] == 63113 && 
b[63114] == 63114 && 
b[63115] == 63115 && 
b[63116] == 63116 && 
b[63117] == 63117 && 
b[63118] == 63118 && 
b[63119] == 63119 && 
b[63120] == 63120 && 
b[63121] == 63121 && 
b[63122] == 63122 && 
b[63123] == 63123 && 
b[63124] == 63124 && 
b[63125] == 63125 && 
b[63126] == 63126 && 
b[63127] == 63127 && 
b[63128] == 63128 && 
b[63129] == 63129 && 
b[63130] == 63130 && 
b[63131] == 63131 && 
b[63132] == 63132 && 
b[63133] == 63133 && 
b[63134] == 63134 && 
b[63135] == 63135 && 
b[63136] == 63136 && 
b[63137] == 63137 && 
b[63138] == 63138 && 
b[63139] == 63139 && 
b[63140] == 63140 && 
b[63141] == 63141 && 
b[63142] == 63142 && 
b[63143] == 63143 && 
b[63144] == 63144 && 
b[63145] == 63145 && 
b[63146] == 63146 && 
b[63147] == 63147 && 
b[63148] == 63148 && 
b[63149] == 63149 && 
b[63150] == 63150 && 
b[63151] == 63151 && 
b[63152] == 63152 && 
b[63153] == 63153 && 
b[63154] == 63154 && 
b[63155] == 63155 && 
b[63156] == 63156 && 
b[63157] == 63157 && 
b[63158] == 63158 && 
b[63159] == 63159 && 
b[63160] == 63160 && 
b[63161] == 63161 && 
b[63162] == 63162 && 
b[63163] == 63163 && 
b[63164] == 63164 && 
b[63165] == 63165 && 
b[63166] == 63166 && 
b[63167] == 63167 && 
b[63168] == 63168 && 
b[63169] == 63169 && 
b[63170] == 63170 && 
b[63171] == 63171 && 
b[63172] == 63172 && 
b[63173] == 63173 && 
b[63174] == 63174 && 
b[63175] == 63175 && 
b[63176] == 63176 && 
b[63177] == 63177 && 
b[63178] == 63178 && 
b[63179] == 63179 && 
b[63180] == 63180 && 
b[63181] == 63181 && 
b[63182] == 63182 && 
b[63183] == 63183 && 
b[63184] == 63184 && 
b[63185] == 63185 && 
b[63186] == 63186 && 
b[63187] == 63187 && 
b[63188] == 63188 && 
b[63189] == 63189 && 
b[63190] == 63190 && 
b[63191] == 63191 && 
b[63192] == 63192 && 
b[63193] == 63193 && 
b[63194] == 63194 && 
b[63195] == 63195 && 
b[63196] == 63196 && 
b[63197] == 63197 && 
b[63198] == 63198 && 
b[63199] == 63199 && 
b[63200] == 63200 && 
b[63201] == 63201 && 
b[63202] == 63202 && 
b[63203] == 63203 && 
b[63204] == 63204 && 
b[63205] == 63205 && 
b[63206] == 63206 && 
b[63207] == 63207 && 
b[63208] == 63208 && 
b[63209] == 63209 && 
b[63210] == 63210 && 
b[63211] == 63211 && 
b[63212] == 63212 && 
b[63213] == 63213 && 
b[63214] == 63214 && 
b[63215] == 63215 && 
b[63216] == 63216 && 
b[63217] == 63217 && 
b[63218] == 63218 && 
b[63219] == 63219 && 
b[63220] == 63220 && 
b[63221] == 63221 && 
b[63222] == 63222 && 
b[63223] == 63223 && 
b[63224] == 63224 && 
b[63225] == 63225 && 
b[63226] == 63226 && 
b[63227] == 63227 && 
b[63228] == 63228 && 
b[63229] == 63229 && 
b[63230] == 63230 && 
b[63231] == 63231 && 
b[63232] == 63232 && 
b[63233] == 63233 && 
b[63234] == 63234 && 
b[63235] == 63235 && 
b[63236] == 63236 && 
b[63237] == 63237 && 
b[63238] == 63238 && 
b[63239] == 63239 && 
b[63240] == 63240 && 
b[63241] == 63241 && 
b[63242] == 63242 && 
b[63243] == 63243 && 
b[63244] == 63244 && 
b[63245] == 63245 && 
b[63246] == 63246 && 
b[63247] == 63247 && 
b[63248] == 63248 && 
b[63249] == 63249 && 
b[63250] == 63250 && 
b[63251] == 63251 && 
b[63252] == 63252 && 
b[63253] == 63253 && 
b[63254] == 63254 && 
b[63255] == 63255 && 
b[63256] == 63256 && 
b[63257] == 63257 && 
b[63258] == 63258 && 
b[63259] == 63259 && 
b[63260] == 63260 && 
b[63261] == 63261 && 
b[63262] == 63262 && 
b[63263] == 63263 && 
b[63264] == 63264 && 
b[63265] == 63265 && 
b[63266] == 63266 && 
b[63267] == 63267 && 
b[63268] == 63268 && 
b[63269] == 63269 && 
b[63270] == 63270 && 
b[63271] == 63271 && 
b[63272] == 63272 && 
b[63273] == 63273 && 
b[63274] == 63274 && 
b[63275] == 63275 && 
b[63276] == 63276 && 
b[63277] == 63277 && 
b[63278] == 63278 && 
b[63279] == 63279 && 
b[63280] == 63280 && 
b[63281] == 63281 && 
b[63282] == 63282 && 
b[63283] == 63283 && 
b[63284] == 63284 && 
b[63285] == 63285 && 
b[63286] == 63286 && 
b[63287] == 63287 && 
b[63288] == 63288 && 
b[63289] == 63289 && 
b[63290] == 63290 && 
b[63291] == 63291 && 
b[63292] == 63292 && 
b[63293] == 63293 && 
b[63294] == 63294 && 
b[63295] == 63295 && 
b[63296] == 63296 && 
b[63297] == 63297 && 
b[63298] == 63298 && 
b[63299] == 63299 && 
b[63300] == 63300 && 
b[63301] == 63301 && 
b[63302] == 63302 && 
b[63303] == 63303 && 
b[63304] == 63304 && 
b[63305] == 63305 && 
b[63306] == 63306 && 
b[63307] == 63307 && 
b[63308] == 63308 && 
b[63309] == 63309 && 
b[63310] == 63310 && 
b[63311] == 63311 && 
b[63312] == 63312 && 
b[63313] == 63313 && 
b[63314] == 63314 && 
b[63315] == 63315 && 
b[63316] == 63316 && 
b[63317] == 63317 && 
b[63318] == 63318 && 
b[63319] == 63319 && 
b[63320] == 63320 && 
b[63321] == 63321 && 
b[63322] == 63322 && 
b[63323] == 63323 && 
b[63324] == 63324 && 
b[63325] == 63325 && 
b[63326] == 63326 && 
b[63327] == 63327 && 
b[63328] == 63328 && 
b[63329] == 63329 && 
b[63330] == 63330 && 
b[63331] == 63331 && 
b[63332] == 63332 && 
b[63333] == 63333 && 
b[63334] == 63334 && 
b[63335] == 63335 && 
b[63336] == 63336 && 
b[63337] == 63337 && 
b[63338] == 63338 && 
b[63339] == 63339 && 
b[63340] == 63340 && 
b[63341] == 63341 && 
b[63342] == 63342 && 
b[63343] == 63343 && 
b[63344] == 63344 && 
b[63345] == 63345 && 
b[63346] == 63346 && 
b[63347] == 63347 && 
b[63348] == 63348 && 
b[63349] == 63349 && 
b[63350] == 63350 && 
b[63351] == 63351 && 
b[63352] == 63352 && 
b[63353] == 63353 && 
b[63354] == 63354 && 
b[63355] == 63355 && 
b[63356] == 63356 && 
b[63357] == 63357 && 
b[63358] == 63358 && 
b[63359] == 63359 && 
b[63360] == 63360 && 
b[63361] == 63361 && 
b[63362] == 63362 && 
b[63363] == 63363 && 
b[63364] == 63364 && 
b[63365] == 63365 && 
b[63366] == 63366 && 
b[63367] == 63367 && 
b[63368] == 63368 && 
b[63369] == 63369 && 
b[63370] == 63370 && 
b[63371] == 63371 && 
b[63372] == 63372 && 
b[63373] == 63373 && 
b[63374] == 63374 && 
b[63375] == 63375 && 
b[63376] == 63376 && 
b[63377] == 63377 && 
b[63378] == 63378 && 
b[63379] == 63379 && 
b[63380] == 63380 && 
b[63381] == 63381 && 
b[63382] == 63382 && 
b[63383] == 63383 && 
b[63384] == 63384 && 
b[63385] == 63385 && 
b[63386] == 63386 && 
b[63387] == 63387 && 
b[63388] == 63388 && 
b[63389] == 63389 && 
b[63390] == 63390 && 
b[63391] == 63391 && 
b[63392] == 63392 && 
b[63393] == 63393 && 
b[63394] == 63394 && 
b[63395] == 63395 && 
b[63396] == 63396 && 
b[63397] == 63397 && 
b[63398] == 63398 && 
b[63399] == 63399 && 
b[63400] == 63400 && 
b[63401] == 63401 && 
b[63402] == 63402 && 
b[63403] == 63403 && 
b[63404] == 63404 && 
b[63405] == 63405 && 
b[63406] == 63406 && 
b[63407] == 63407 && 
b[63408] == 63408 && 
b[63409] == 63409 && 
b[63410] == 63410 && 
b[63411] == 63411 && 
b[63412] == 63412 && 
b[63413] == 63413 && 
b[63414] == 63414 && 
b[63415] == 63415 && 
b[63416] == 63416 && 
b[63417] == 63417 && 
b[63418] == 63418 && 
b[63419] == 63419 && 
b[63420] == 63420 && 
b[63421] == 63421 && 
b[63422] == 63422 && 
b[63423] == 63423 && 
b[63424] == 63424 && 
b[63425] == 63425 && 
b[63426] == 63426 && 
b[63427] == 63427 && 
b[63428] == 63428 && 
b[63429] == 63429 && 
b[63430] == 63430 && 
b[63431] == 63431 && 
b[63432] == 63432 && 
b[63433] == 63433 && 
b[63434] == 63434 && 
b[63435] == 63435 && 
b[63436] == 63436 && 
b[63437] == 63437 && 
b[63438] == 63438 && 
b[63439] == 63439 && 
b[63440] == 63440 && 
b[63441] == 63441 && 
b[63442] == 63442 && 
b[63443] == 63443 && 
b[63444] == 63444 && 
b[63445] == 63445 && 
b[63446] == 63446 && 
b[63447] == 63447 && 
b[63448] == 63448 && 
b[63449] == 63449 && 
b[63450] == 63450 && 
b[63451] == 63451 && 
b[63452] == 63452 && 
b[63453] == 63453 && 
b[63454] == 63454 && 
b[63455] == 63455 && 
b[63456] == 63456 && 
b[63457] == 63457 && 
b[63458] == 63458 && 
b[63459] == 63459 && 
b[63460] == 63460 && 
b[63461] == 63461 && 
b[63462] == 63462 && 
b[63463] == 63463 && 
b[63464] == 63464 && 
b[63465] == 63465 && 
b[63466] == 63466 && 
b[63467] == 63467 && 
b[63468] == 63468 && 
b[63469] == 63469 && 
b[63470] == 63470 && 
b[63471] == 63471 && 
b[63472] == 63472 && 
b[63473] == 63473 && 
b[63474] == 63474 && 
b[63475] == 63475 && 
b[63476] == 63476 && 
b[63477] == 63477 && 
b[63478] == 63478 && 
b[63479] == 63479 && 
b[63480] == 63480 && 
b[63481] == 63481 && 
b[63482] == 63482 && 
b[63483] == 63483 && 
b[63484] == 63484 && 
b[63485] == 63485 && 
b[63486] == 63486 && 
b[63487] == 63487 && 
b[63488] == 63488 && 
b[63489] == 63489 && 
b[63490] == 63490 && 
b[63491] == 63491 && 
b[63492] == 63492 && 
b[63493] == 63493 && 
b[63494] == 63494 && 
b[63495] == 63495 && 
b[63496] == 63496 && 
b[63497] == 63497 && 
b[63498] == 63498 && 
b[63499] == 63499 && 
b[63500] == 63500 && 
b[63501] == 63501 && 
b[63502] == 63502 && 
b[63503] == 63503 && 
b[63504] == 63504 && 
b[63505] == 63505 && 
b[63506] == 63506 && 
b[63507] == 63507 && 
b[63508] == 63508 && 
b[63509] == 63509 && 
b[63510] == 63510 && 
b[63511] == 63511 && 
b[63512] == 63512 && 
b[63513] == 63513 && 
b[63514] == 63514 && 
b[63515] == 63515 && 
b[63516] == 63516 && 
b[63517] == 63517 && 
b[63518] == 63518 && 
b[63519] == 63519 && 
b[63520] == 63520 && 
b[63521] == 63521 && 
b[63522] == 63522 && 
b[63523] == 63523 && 
b[63524] == 63524 && 
b[63525] == 63525 && 
b[63526] == 63526 && 
b[63527] == 63527 && 
b[63528] == 63528 && 
b[63529] == 63529 && 
b[63530] == 63530 && 
b[63531] == 63531 && 
b[63532] == 63532 && 
b[63533] == 63533 && 
b[63534] == 63534 && 
b[63535] == 63535 && 
b[63536] == 63536 && 
b[63537] == 63537 && 
b[63538] == 63538 && 
b[63539] == 63539 && 
b[63540] == 63540 && 
b[63541] == 63541 && 
b[63542] == 63542 && 
b[63543] == 63543 && 
b[63544] == 63544 && 
b[63545] == 63545 && 
b[63546] == 63546 && 
b[63547] == 63547 && 
b[63548] == 63548 && 
b[63549] == 63549 && 
b[63550] == 63550 && 
b[63551] == 63551 && 
b[63552] == 63552 && 
b[63553] == 63553 && 
b[63554] == 63554 && 
b[63555] == 63555 && 
b[63556] == 63556 && 
b[63557] == 63557 && 
b[63558] == 63558 && 
b[63559] == 63559 && 
b[63560] == 63560 && 
b[63561] == 63561 && 
b[63562] == 63562 && 
b[63563] == 63563 && 
b[63564] == 63564 && 
b[63565] == 63565 && 
b[63566] == 63566 && 
b[63567] == 63567 && 
b[63568] == 63568 && 
b[63569] == 63569 && 
b[63570] == 63570 && 
b[63571] == 63571 && 
b[63572] == 63572 && 
b[63573] == 63573 && 
b[63574] == 63574 && 
b[63575] == 63575 && 
b[63576] == 63576 && 
b[63577] == 63577 && 
b[63578] == 63578 && 
b[63579] == 63579 && 
b[63580] == 63580 && 
b[63581] == 63581 && 
b[63582] == 63582 && 
b[63583] == 63583 && 
b[63584] == 63584 && 
b[63585] == 63585 && 
b[63586] == 63586 && 
b[63587] == 63587 && 
b[63588] == 63588 && 
b[63589] == 63589 && 
b[63590] == 63590 && 
b[63591] == 63591 && 
b[63592] == 63592 && 
b[63593] == 63593 && 
b[63594] == 63594 && 
b[63595] == 63595 && 
b[63596] == 63596 && 
b[63597] == 63597 && 
b[63598] == 63598 && 
b[63599] == 63599 && 
b[63600] == 63600 && 
b[63601] == 63601 && 
b[63602] == 63602 && 
b[63603] == 63603 && 
b[63604] == 63604 && 
b[63605] == 63605 && 
b[63606] == 63606 && 
b[63607] == 63607 && 
b[63608] == 63608 && 
b[63609] == 63609 && 
b[63610] == 63610 && 
b[63611] == 63611 && 
b[63612] == 63612 && 
b[63613] == 63613 && 
b[63614] == 63614 && 
b[63615] == 63615 && 
b[63616] == 63616 && 
b[63617] == 63617 && 
b[63618] == 63618 && 
b[63619] == 63619 && 
b[63620] == 63620 && 
b[63621] == 63621 && 
b[63622] == 63622 && 
b[63623] == 63623 && 
b[63624] == 63624 && 
b[63625] == 63625 && 
b[63626] == 63626 && 
b[63627] == 63627 && 
b[63628] == 63628 && 
b[63629] == 63629 && 
b[63630] == 63630 && 
b[63631] == 63631 && 
b[63632] == 63632 && 
b[63633] == 63633 && 
b[63634] == 63634 && 
b[63635] == 63635 && 
b[63636] == 63636 && 
b[63637] == 63637 && 
b[63638] == 63638 && 
b[63639] == 63639 && 
b[63640] == 63640 && 
b[63641] == 63641 && 
b[63642] == 63642 && 
b[63643] == 63643 && 
b[63644] == 63644 && 
b[63645] == 63645 && 
b[63646] == 63646 && 
b[63647] == 63647 && 
b[63648] == 63648 && 
b[63649] == 63649 && 
b[63650] == 63650 && 
b[63651] == 63651 && 
b[63652] == 63652 && 
b[63653] == 63653 && 
b[63654] == 63654 && 
b[63655] == 63655 && 
b[63656] == 63656 && 
b[63657] == 63657 && 
b[63658] == 63658 && 
b[63659] == 63659 && 
b[63660] == 63660 && 
b[63661] == 63661 && 
b[63662] == 63662 && 
b[63663] == 63663 && 
b[63664] == 63664 && 
b[63665] == 63665 && 
b[63666] == 63666 && 
b[63667] == 63667 && 
b[63668] == 63668 && 
b[63669] == 63669 && 
b[63670] == 63670 && 
b[63671] == 63671 && 
b[63672] == 63672 && 
b[63673] == 63673 && 
b[63674] == 63674 && 
b[63675] == 63675 && 
b[63676] == 63676 && 
b[63677] == 63677 && 
b[63678] == 63678 && 
b[63679] == 63679 && 
b[63680] == 63680 && 
b[63681] == 63681 && 
b[63682] == 63682 && 
b[63683] == 63683 && 
b[63684] == 63684 && 
b[63685] == 63685 && 
b[63686] == 63686 && 
b[63687] == 63687 && 
b[63688] == 63688 && 
b[63689] == 63689 && 
b[63690] == 63690 && 
b[63691] == 63691 && 
b[63692] == 63692 && 
b[63693] == 63693 && 
b[63694] == 63694 && 
b[63695] == 63695 && 
b[63696] == 63696 && 
b[63697] == 63697 && 
b[63698] == 63698 && 
b[63699] == 63699 && 
b[63700] == 63700 && 
b[63701] == 63701 && 
b[63702] == 63702 && 
b[63703] == 63703 && 
b[63704] == 63704 && 
b[63705] == 63705 && 
b[63706] == 63706 && 
b[63707] == 63707 && 
b[63708] == 63708 && 
b[63709] == 63709 && 
b[63710] == 63710 && 
b[63711] == 63711 && 
b[63712] == 63712 && 
b[63713] == 63713 && 
b[63714] == 63714 && 
b[63715] == 63715 && 
b[63716] == 63716 && 
b[63717] == 63717 && 
b[63718] == 63718 && 
b[63719] == 63719 && 
b[63720] == 63720 && 
b[63721] == 63721 && 
b[63722] == 63722 && 
b[63723] == 63723 && 
b[63724] == 63724 && 
b[63725] == 63725 && 
b[63726] == 63726 && 
b[63727] == 63727 && 
b[63728] == 63728 && 
b[63729] == 63729 && 
b[63730] == 63730 && 
b[63731] == 63731 && 
b[63732] == 63732 && 
b[63733] == 63733 && 
b[63734] == 63734 && 
b[63735] == 63735 && 
b[63736] == 63736 && 
b[63737] == 63737 && 
b[63738] == 63738 && 
b[63739] == 63739 && 
b[63740] == 63740 && 
b[63741] == 63741 && 
b[63742] == 63742 && 
b[63743] == 63743 && 
b[63744] == 63744 && 
b[63745] == 63745 && 
b[63746] == 63746 && 
b[63747] == 63747 && 
b[63748] == 63748 && 
b[63749] == 63749 && 
b[63750] == 63750 && 
b[63751] == 63751 && 
b[63752] == 63752 && 
b[63753] == 63753 && 
b[63754] == 63754 && 
b[63755] == 63755 && 
b[63756] == 63756 && 
b[63757] == 63757 && 
b[63758] == 63758 && 
b[63759] == 63759 && 
b[63760] == 63760 && 
b[63761] == 63761 && 
b[63762] == 63762 && 
b[63763] == 63763 && 
b[63764] == 63764 && 
b[63765] == 63765 && 
b[63766] == 63766 && 
b[63767] == 63767 && 
b[63768] == 63768 && 
b[63769] == 63769 && 
b[63770] == 63770 && 
b[63771] == 63771 && 
b[63772] == 63772 && 
b[63773] == 63773 && 
b[63774] == 63774 && 
b[63775] == 63775 && 
b[63776] == 63776 && 
b[63777] == 63777 && 
b[63778] == 63778 && 
b[63779] == 63779 && 
b[63780] == 63780 && 
b[63781] == 63781 && 
b[63782] == 63782 && 
b[63783] == 63783 && 
b[63784] == 63784 && 
b[63785] == 63785 && 
b[63786] == 63786 && 
b[63787] == 63787 && 
b[63788] == 63788 && 
b[63789] == 63789 && 
b[63790] == 63790 && 
b[63791] == 63791 && 
b[63792] == 63792 && 
b[63793] == 63793 && 
b[63794] == 63794 && 
b[63795] == 63795 && 
b[63796] == 63796 && 
b[63797] == 63797 && 
b[63798] == 63798 && 
b[63799] == 63799 && 
b[63800] == 63800 && 
b[63801] == 63801 && 
b[63802] == 63802 && 
b[63803] == 63803 && 
b[63804] == 63804 && 
b[63805] == 63805 && 
b[63806] == 63806 && 
b[63807] == 63807 && 
b[63808] == 63808 && 
b[63809] == 63809 && 
b[63810] == 63810 && 
b[63811] == 63811 && 
b[63812] == 63812 && 
b[63813] == 63813 && 
b[63814] == 63814 && 
b[63815] == 63815 && 
b[63816] == 63816 && 
b[63817] == 63817 && 
b[63818] == 63818 && 
b[63819] == 63819 && 
b[63820] == 63820 && 
b[63821] == 63821 && 
b[63822] == 63822 && 
b[63823] == 63823 && 
b[63824] == 63824 && 
b[63825] == 63825 && 
b[63826] == 63826 && 
b[63827] == 63827 && 
b[63828] == 63828 && 
b[63829] == 63829 && 
b[63830] == 63830 && 
b[63831] == 63831 && 
b[63832] == 63832 && 
b[63833] == 63833 && 
b[63834] == 63834 && 
b[63835] == 63835 && 
b[63836] == 63836 && 
b[63837] == 63837 && 
b[63838] == 63838 && 
b[63839] == 63839 && 
b[63840] == 63840 && 
b[63841] == 63841 && 
b[63842] == 63842 && 
b[63843] == 63843 && 
b[63844] == 63844 && 
b[63845] == 63845 && 
b[63846] == 63846 && 
b[63847] == 63847 && 
b[63848] == 63848 && 
b[63849] == 63849 && 
b[63850] == 63850 && 
b[63851] == 63851 && 
b[63852] == 63852 && 
b[63853] == 63853 && 
b[63854] == 63854 && 
b[63855] == 63855 && 
b[63856] == 63856 && 
b[63857] == 63857 && 
b[63858] == 63858 && 
b[63859] == 63859 && 
b[63860] == 63860 && 
b[63861] == 63861 && 
b[63862] == 63862 && 
b[63863] == 63863 && 
b[63864] == 63864 && 
b[63865] == 63865 && 
b[63866] == 63866 && 
b[63867] == 63867 && 
b[63868] == 63868 && 
b[63869] == 63869 && 
b[63870] == 63870 && 
b[63871] == 63871 && 
b[63872] == 63872 && 
b[63873] == 63873 && 
b[63874] == 63874 && 
b[63875] == 63875 && 
b[63876] == 63876 && 
b[63877] == 63877 && 
b[63878] == 63878 && 
b[63879] == 63879 && 
b[63880] == 63880 && 
b[63881] == 63881 && 
b[63882] == 63882 && 
b[63883] == 63883 && 
b[63884] == 63884 && 
b[63885] == 63885 && 
b[63886] == 63886 && 
b[63887] == 63887 && 
b[63888] == 63888 && 
b[63889] == 63889 && 
b[63890] == 63890 && 
b[63891] == 63891 && 
b[63892] == 63892 && 
b[63893] == 63893 && 
b[63894] == 63894 && 
b[63895] == 63895 && 
b[63896] == 63896 && 
b[63897] == 63897 && 
b[63898] == 63898 && 
b[63899] == 63899 && 
b[63900] == 63900 && 
b[63901] == 63901 && 
b[63902] == 63902 && 
b[63903] == 63903 && 
b[63904] == 63904 && 
b[63905] == 63905 && 
b[63906] == 63906 && 
b[63907] == 63907 && 
b[63908] == 63908 && 
b[63909] == 63909 && 
b[63910] == 63910 && 
b[63911] == 63911 && 
b[63912] == 63912 && 
b[63913] == 63913 && 
b[63914] == 63914 && 
b[63915] == 63915 && 
b[63916] == 63916 && 
b[63917] == 63917 && 
b[63918] == 63918 && 
b[63919] == 63919 && 
b[63920] == 63920 && 
b[63921] == 63921 && 
b[63922] == 63922 && 
b[63923] == 63923 && 
b[63924] == 63924 && 
b[63925] == 63925 && 
b[63926] == 63926 && 
b[63927] == 63927 && 
b[63928] == 63928 && 
b[63929] == 63929 && 
b[63930] == 63930 && 
b[63931] == 63931 && 
b[63932] == 63932 && 
b[63933] == 63933 && 
b[63934] == 63934 && 
b[63935] == 63935 && 
b[63936] == 63936 && 
b[63937] == 63937 && 
b[63938] == 63938 && 
b[63939] == 63939 && 
b[63940] == 63940 && 
b[63941] == 63941 && 
b[63942] == 63942 && 
b[63943] == 63943 && 
b[63944] == 63944 && 
b[63945] == 63945 && 
b[63946] == 63946 && 
b[63947] == 63947 && 
b[63948] == 63948 && 
b[63949] == 63949 && 
b[63950] == 63950 && 
b[63951] == 63951 && 
b[63952] == 63952 && 
b[63953] == 63953 && 
b[63954] == 63954 && 
b[63955] == 63955 && 
b[63956] == 63956 && 
b[63957] == 63957 && 
b[63958] == 63958 && 
b[63959] == 63959 && 
b[63960] == 63960 && 
b[63961] == 63961 && 
b[63962] == 63962 && 
b[63963] == 63963 && 
b[63964] == 63964 && 
b[63965] == 63965 && 
b[63966] == 63966 && 
b[63967] == 63967 && 
b[63968] == 63968 && 
b[63969] == 63969 && 
b[63970] == 63970 && 
b[63971] == 63971 && 
b[63972] == 63972 && 
b[63973] == 63973 && 
b[63974] == 63974 && 
b[63975] == 63975 && 
b[63976] == 63976 && 
b[63977] == 63977 && 
b[63978] == 63978 && 
b[63979] == 63979 && 
b[63980] == 63980 && 
b[63981] == 63981 && 
b[63982] == 63982 && 
b[63983] == 63983 && 
b[63984] == 63984 && 
b[63985] == 63985 && 
b[63986] == 63986 && 
b[63987] == 63987 && 
b[63988] == 63988 && 
b[63989] == 63989 && 
b[63990] == 63990 && 
b[63991] == 63991 && 
b[63992] == 63992 && 
b[63993] == 63993 && 
b[63994] == 63994 && 
b[63995] == 63995 && 
b[63996] == 63996 && 
b[63997] == 63997 && 
b[63998] == 63998 && 
b[63999] == 63999 && 
b[64000] == 64000 && 
b[64001] == 64001 && 
b[64002] == 64002 && 
b[64003] == 64003 && 
b[64004] == 64004 && 
b[64005] == 64005 && 
b[64006] == 64006 && 
b[64007] == 64007 && 
b[64008] == 64008 && 
b[64009] == 64009 && 
b[64010] == 64010 && 
b[64011] == 64011 && 
b[64012] == 64012 && 
b[64013] == 64013 && 
b[64014] == 64014 && 
b[64015] == 64015 && 
b[64016] == 64016 && 
b[64017] == 64017 && 
b[64018] == 64018 && 
b[64019] == 64019 && 
b[64020] == 64020 && 
b[64021] == 64021 && 
b[64022] == 64022 && 
b[64023] == 64023 && 
b[64024] == 64024 && 
b[64025] == 64025 && 
b[64026] == 64026 && 
b[64027] == 64027 && 
b[64028] == 64028 && 
b[64029] == 64029 && 
b[64030] == 64030 && 
b[64031] == 64031 && 
b[64032] == 64032 && 
b[64033] == 64033 && 
b[64034] == 64034 && 
b[64035] == 64035 && 
b[64036] == 64036 && 
b[64037] == 64037 && 
b[64038] == 64038 && 
b[64039] == 64039 && 
b[64040] == 64040 && 
b[64041] == 64041 && 
b[64042] == 64042 && 
b[64043] == 64043 && 
b[64044] == 64044 && 
b[64045] == 64045 && 
b[64046] == 64046 && 
b[64047] == 64047 && 
b[64048] == 64048 && 
b[64049] == 64049 && 
b[64050] == 64050 && 
b[64051] == 64051 && 
b[64052] == 64052 && 
b[64053] == 64053 && 
b[64054] == 64054 && 
b[64055] == 64055 && 
b[64056] == 64056 && 
b[64057] == 64057 && 
b[64058] == 64058 && 
b[64059] == 64059 && 
b[64060] == 64060 && 
b[64061] == 64061 && 
b[64062] == 64062 && 
b[64063] == 64063 && 
b[64064] == 64064 && 
b[64065] == 64065 && 
b[64066] == 64066 && 
b[64067] == 64067 && 
b[64068] == 64068 && 
b[64069] == 64069 && 
b[64070] == 64070 && 
b[64071] == 64071 && 
b[64072] == 64072 && 
b[64073] == 64073 && 
b[64074] == 64074 && 
b[64075] == 64075 && 
b[64076] == 64076 && 
b[64077] == 64077 && 
b[64078] == 64078 && 
b[64079] == 64079 && 
b[64080] == 64080 && 
b[64081] == 64081 && 
b[64082] == 64082 && 
b[64083] == 64083 && 
b[64084] == 64084 && 
b[64085] == 64085 && 
b[64086] == 64086 && 
b[64087] == 64087 && 
b[64088] == 64088 && 
b[64089] == 64089 && 
b[64090] == 64090 && 
b[64091] == 64091 && 
b[64092] == 64092 && 
b[64093] == 64093 && 
b[64094] == 64094 && 
b[64095] == 64095 && 
b[64096] == 64096 && 
b[64097] == 64097 && 
b[64098] == 64098 && 
b[64099] == 64099 && 
b[64100] == 64100 && 
b[64101] == 64101 && 
b[64102] == 64102 && 
b[64103] == 64103 && 
b[64104] == 64104 && 
b[64105] == 64105 && 
b[64106] == 64106 && 
b[64107] == 64107 && 
b[64108] == 64108 && 
b[64109] == 64109 && 
b[64110] == 64110 && 
b[64111] == 64111 && 
b[64112] == 64112 && 
b[64113] == 64113 && 
b[64114] == 64114 && 
b[64115] == 64115 && 
b[64116] == 64116 && 
b[64117] == 64117 && 
b[64118] == 64118 && 
b[64119] == 64119 && 
b[64120] == 64120 && 
b[64121] == 64121 && 
b[64122] == 64122 && 
b[64123] == 64123 && 
b[64124] == 64124 && 
b[64125] == 64125 && 
b[64126] == 64126 && 
b[64127] == 64127 && 
b[64128] == 64128 && 
b[64129] == 64129 && 
b[64130] == 64130 && 
b[64131] == 64131 && 
b[64132] == 64132 && 
b[64133] == 64133 && 
b[64134] == 64134 && 
b[64135] == 64135 && 
b[64136] == 64136 && 
b[64137] == 64137 && 
b[64138] == 64138 && 
b[64139] == 64139 && 
b[64140] == 64140 && 
b[64141] == 64141 && 
b[64142] == 64142 && 
b[64143] == 64143 && 
b[64144] == 64144 && 
b[64145] == 64145 && 
b[64146] == 64146 && 
b[64147] == 64147 && 
b[64148] == 64148 && 
b[64149] == 64149 && 
b[64150] == 64150 && 
b[64151] == 64151 && 
b[64152] == 64152 && 
b[64153] == 64153 && 
b[64154] == 64154 && 
b[64155] == 64155 && 
b[64156] == 64156 && 
b[64157] == 64157 && 
b[64158] == 64158 && 
b[64159] == 64159 && 
b[64160] == 64160 && 
b[64161] == 64161 && 
b[64162] == 64162 && 
b[64163] == 64163 && 
b[64164] == 64164 && 
b[64165] == 64165 && 
b[64166] == 64166 && 
b[64167] == 64167 && 
b[64168] == 64168 && 
b[64169] == 64169 && 
b[64170] == 64170 && 
b[64171] == 64171 && 
b[64172] == 64172 && 
b[64173] == 64173 && 
b[64174] == 64174 && 
b[64175] == 64175 && 
b[64176] == 64176 && 
b[64177] == 64177 && 
b[64178] == 64178 && 
b[64179] == 64179 && 
b[64180] == 64180 && 
b[64181] == 64181 && 
b[64182] == 64182 && 
b[64183] == 64183 && 
b[64184] == 64184 && 
b[64185] == 64185 && 
b[64186] == 64186 && 
b[64187] == 64187 && 
b[64188] == 64188 && 
b[64189] == 64189 && 
b[64190] == 64190 && 
b[64191] == 64191 && 
b[64192] == 64192 && 
b[64193] == 64193 && 
b[64194] == 64194 && 
b[64195] == 64195 && 
b[64196] == 64196 && 
b[64197] == 64197 && 
b[64198] == 64198 && 
b[64199] == 64199 && 
b[64200] == 64200 && 
b[64201] == 64201 && 
b[64202] == 64202 && 
b[64203] == 64203 && 
b[64204] == 64204 && 
b[64205] == 64205 && 
b[64206] == 64206 && 
b[64207] == 64207 && 
b[64208] == 64208 && 
b[64209] == 64209 && 
b[64210] == 64210 && 
b[64211] == 64211 && 
b[64212] == 64212 && 
b[64213] == 64213 && 
b[64214] == 64214 && 
b[64215] == 64215 && 
b[64216] == 64216 && 
b[64217] == 64217 && 
b[64218] == 64218 && 
b[64219] == 64219 && 
b[64220] == 64220 && 
b[64221] == 64221 && 
b[64222] == 64222 && 
b[64223] == 64223 && 
b[64224] == 64224 && 
b[64225] == 64225 && 
b[64226] == 64226 && 
b[64227] == 64227 && 
b[64228] == 64228 && 
b[64229] == 64229 && 
b[64230] == 64230 && 
b[64231] == 64231 && 
b[64232] == 64232 && 
b[64233] == 64233 && 
b[64234] == 64234 && 
b[64235] == 64235 && 
b[64236] == 64236 && 
b[64237] == 64237 && 
b[64238] == 64238 && 
b[64239] == 64239 && 
b[64240] == 64240 && 
b[64241] == 64241 && 
b[64242] == 64242 && 
b[64243] == 64243 && 
b[64244] == 64244 && 
b[64245] == 64245 && 
b[64246] == 64246 && 
b[64247] == 64247 && 
b[64248] == 64248 && 
b[64249] == 64249 && 
b[64250] == 64250 && 
b[64251] == 64251 && 
b[64252] == 64252 && 
b[64253] == 64253 && 
b[64254] == 64254 && 
b[64255] == 64255 && 
b[64256] == 64256 && 
b[64257] == 64257 && 
b[64258] == 64258 && 
b[64259] == 64259 && 
b[64260] == 64260 && 
b[64261] == 64261 && 
b[64262] == 64262 && 
b[64263] == 64263 && 
b[64264] == 64264 && 
b[64265] == 64265 && 
b[64266] == 64266 && 
b[64267] == 64267 && 
b[64268] == 64268 && 
b[64269] == 64269 && 
b[64270] == 64270 && 
b[64271] == 64271 && 
b[64272] == 64272 && 
b[64273] == 64273 && 
b[64274] == 64274 && 
b[64275] == 64275 && 
b[64276] == 64276 && 
b[64277] == 64277 && 
b[64278] == 64278 && 
b[64279] == 64279 && 
b[64280] == 64280 && 
b[64281] == 64281 && 
b[64282] == 64282 && 
b[64283] == 64283 && 
b[64284] == 64284 && 
b[64285] == 64285 && 
b[64286] == 64286 && 
b[64287] == 64287 && 
b[64288] == 64288 && 
b[64289] == 64289 && 
b[64290] == 64290 && 
b[64291] == 64291 && 
b[64292] == 64292 && 
b[64293] == 64293 && 
b[64294] == 64294 && 
b[64295] == 64295 && 
b[64296] == 64296 && 
b[64297] == 64297 && 
b[64298] == 64298 && 
b[64299] == 64299 && 
b[64300] == 64300 && 
b[64301] == 64301 && 
b[64302] == 64302 && 
b[64303] == 64303 && 
b[64304] == 64304 && 
b[64305] == 64305 && 
b[64306] == 64306 && 
b[64307] == 64307 && 
b[64308] == 64308 && 
b[64309] == 64309 && 
b[64310] == 64310 && 
b[64311] == 64311 && 
b[64312] == 64312 && 
b[64313] == 64313 && 
b[64314] == 64314 && 
b[64315] == 64315 && 
b[64316] == 64316 && 
b[64317] == 64317 && 
b[64318] == 64318 && 
b[64319] == 64319 && 
b[64320] == 64320 && 
b[64321] == 64321 && 
b[64322] == 64322 && 
b[64323] == 64323 && 
b[64324] == 64324 && 
b[64325] == 64325 && 
b[64326] == 64326 && 
b[64327] == 64327 && 
b[64328] == 64328 && 
b[64329] == 64329 && 
b[64330] == 64330 && 
b[64331] == 64331 && 
b[64332] == 64332 && 
b[64333] == 64333 && 
b[64334] == 64334 && 
b[64335] == 64335 && 
b[64336] == 64336 && 
b[64337] == 64337 && 
b[64338] == 64338 && 
b[64339] == 64339 && 
b[64340] == 64340 && 
b[64341] == 64341 && 
b[64342] == 64342 && 
b[64343] == 64343 && 
b[64344] == 64344 && 
b[64345] == 64345 && 
b[64346] == 64346 && 
b[64347] == 64347 && 
b[64348] == 64348 && 
b[64349] == 64349 && 
b[64350] == 64350 && 
b[64351] == 64351 && 
b[64352] == 64352 && 
b[64353] == 64353 && 
b[64354] == 64354 && 
b[64355] == 64355 && 
b[64356] == 64356 && 
b[64357] == 64357 && 
b[64358] == 64358 && 
b[64359] == 64359 && 
b[64360] == 64360 && 
b[64361] == 64361 && 
b[64362] == 64362 && 
b[64363] == 64363 && 
b[64364] == 64364 && 
b[64365] == 64365 && 
b[64366] == 64366 && 
b[64367] == 64367 && 
b[64368] == 64368 && 
b[64369] == 64369 && 
b[64370] == 64370 && 
b[64371] == 64371 && 
b[64372] == 64372 && 
b[64373] == 64373 && 
b[64374] == 64374 && 
b[64375] == 64375 && 
b[64376] == 64376 && 
b[64377] == 64377 && 
b[64378] == 64378 && 
b[64379] == 64379 && 
b[64380] == 64380 && 
b[64381] == 64381 && 
b[64382] == 64382 && 
b[64383] == 64383 && 
b[64384] == 64384 && 
b[64385] == 64385 && 
b[64386] == 64386 && 
b[64387] == 64387 && 
b[64388] == 64388 && 
b[64389] == 64389 && 
b[64390] == 64390 && 
b[64391] == 64391 && 
b[64392] == 64392 && 
b[64393] == 64393 && 
b[64394] == 64394 && 
b[64395] == 64395 && 
b[64396] == 64396 && 
b[64397] == 64397 && 
b[64398] == 64398 && 
b[64399] == 64399 && 
b[64400] == 64400 && 
b[64401] == 64401 && 
b[64402] == 64402 && 
b[64403] == 64403 && 
b[64404] == 64404 && 
b[64405] == 64405 && 
b[64406] == 64406 && 
b[64407] == 64407 && 
b[64408] == 64408 && 
b[64409] == 64409 && 
b[64410] == 64410 && 
b[64411] == 64411 && 
b[64412] == 64412 && 
b[64413] == 64413 && 
b[64414] == 64414 && 
b[64415] == 64415 && 
b[64416] == 64416 && 
b[64417] == 64417 && 
b[64418] == 64418 && 
b[64419] == 64419 && 
b[64420] == 64420 && 
b[64421] == 64421 && 
b[64422] == 64422 && 
b[64423] == 64423 && 
b[64424] == 64424 && 
b[64425] == 64425 && 
b[64426] == 64426 && 
b[64427] == 64427 && 
b[64428] == 64428 && 
b[64429] == 64429 && 
b[64430] == 64430 && 
b[64431] == 64431 && 
b[64432] == 64432 && 
b[64433] == 64433 && 
b[64434] == 64434 && 
b[64435] == 64435 && 
b[64436] == 64436 && 
b[64437] == 64437 && 
b[64438] == 64438 && 
b[64439] == 64439 && 
b[64440] == 64440 && 
b[64441] == 64441 && 
b[64442] == 64442 && 
b[64443] == 64443 && 
b[64444] == 64444 && 
b[64445] == 64445 && 
b[64446] == 64446 && 
b[64447] == 64447 && 
b[64448] == 64448 && 
b[64449] == 64449 && 
b[64450] == 64450 && 
b[64451] == 64451 && 
b[64452] == 64452 && 
b[64453] == 64453 && 
b[64454] == 64454 && 
b[64455] == 64455 && 
b[64456] == 64456 && 
b[64457] == 64457 && 
b[64458] == 64458 && 
b[64459] == 64459 && 
b[64460] == 64460 && 
b[64461] == 64461 && 
b[64462] == 64462 && 
b[64463] == 64463 && 
b[64464] == 64464 && 
b[64465] == 64465 && 
b[64466] == 64466 && 
b[64467] == 64467 && 
b[64468] == 64468 && 
b[64469] == 64469 && 
b[64470] == 64470 && 
b[64471] == 64471 && 
b[64472] == 64472 && 
b[64473] == 64473 && 
b[64474] == 64474 && 
b[64475] == 64475 && 
b[64476] == 64476 && 
b[64477] == 64477 && 
b[64478] == 64478 && 
b[64479] == 64479 && 
b[64480] == 64480 && 
b[64481] == 64481 && 
b[64482] == 64482 && 
b[64483] == 64483 && 
b[64484] == 64484 && 
b[64485] == 64485 && 
b[64486] == 64486 && 
b[64487] == 64487 && 
b[64488] == 64488 && 
b[64489] == 64489 && 
b[64490] == 64490 && 
b[64491] == 64491 && 
b[64492] == 64492 && 
b[64493] == 64493 && 
b[64494] == 64494 && 
b[64495] == 64495 && 
b[64496] == 64496 && 
b[64497] == 64497 && 
b[64498] == 64498 && 
b[64499] == 64499 && 
b[64500] == 64500 && 
b[64501] == 64501 && 
b[64502] == 64502 && 
b[64503] == 64503 && 
b[64504] == 64504 && 
b[64505] == 64505 && 
b[64506] == 64506 && 
b[64507] == 64507 && 
b[64508] == 64508 && 
b[64509] == 64509 && 
b[64510] == 64510 && 
b[64511] == 64511 && 
b[64512] == 64512 && 
b[64513] == 64513 && 
b[64514] == 64514 && 
b[64515] == 64515 && 
b[64516] == 64516 && 
b[64517] == 64517 && 
b[64518] == 64518 && 
b[64519] == 64519 && 
b[64520] == 64520 && 
b[64521] == 64521 && 
b[64522] == 64522 && 
b[64523] == 64523 && 
b[64524] == 64524 && 
b[64525] == 64525 && 
b[64526] == 64526 && 
b[64527] == 64527 && 
b[64528] == 64528 && 
b[64529] == 64529 && 
b[64530] == 64530 && 
b[64531] == 64531 && 
b[64532] == 64532 && 
b[64533] == 64533 && 
b[64534] == 64534 && 
b[64535] == 64535 && 
b[64536] == 64536 && 
b[64537] == 64537 && 
b[64538] == 64538 && 
b[64539] == 64539 && 
b[64540] == 64540 && 
b[64541] == 64541 && 
b[64542] == 64542 && 
b[64543] == 64543 && 
b[64544] == 64544 && 
b[64545] == 64545 && 
b[64546] == 64546 && 
b[64547] == 64547 && 
b[64548] == 64548 && 
b[64549] == 64549 && 
b[64550] == 64550 && 
b[64551] == 64551 && 
b[64552] == 64552 && 
b[64553] == 64553 && 
b[64554] == 64554 && 
b[64555] == 64555 && 
b[64556] == 64556 && 
b[64557] == 64557 && 
b[64558] == 64558 && 
b[64559] == 64559 && 
b[64560] == 64560 && 
b[64561] == 64561 && 
b[64562] == 64562 && 
b[64563] == 64563 && 
b[64564] == 64564 && 
b[64565] == 64565 && 
b[64566] == 64566 && 
b[64567] == 64567 && 
b[64568] == 64568 && 
b[64569] == 64569 && 
b[64570] == 64570 && 
b[64571] == 64571 && 
b[64572] == 64572 && 
b[64573] == 64573 && 
b[64574] == 64574 && 
b[64575] == 64575 && 
b[64576] == 64576 && 
b[64577] == 64577 && 
b[64578] == 64578 && 
b[64579] == 64579 && 
b[64580] == 64580 && 
b[64581] == 64581 && 
b[64582] == 64582 && 
b[64583] == 64583 && 
b[64584] == 64584 && 
b[64585] == 64585 && 
b[64586] == 64586 && 
b[64587] == 64587 && 
b[64588] == 64588 && 
b[64589] == 64589 && 
b[64590] == 64590 && 
b[64591] == 64591 && 
b[64592] == 64592 && 
b[64593] == 64593 && 
b[64594] == 64594 && 
b[64595] == 64595 && 
b[64596] == 64596 && 
b[64597] == 64597 && 
b[64598] == 64598 && 
b[64599] == 64599 && 
b[64600] == 64600 && 
b[64601] == 64601 && 
b[64602] == 64602 && 
b[64603] == 64603 && 
b[64604] == 64604 && 
b[64605] == 64605 && 
b[64606] == 64606 && 
b[64607] == 64607 && 
b[64608] == 64608 && 
b[64609] == 64609 && 
b[64610] == 64610 && 
b[64611] == 64611 && 
b[64612] == 64612 && 
b[64613] == 64613 && 
b[64614] == 64614 && 
b[64615] == 64615 && 
b[64616] == 64616 && 
b[64617] == 64617 && 
b[64618] == 64618 && 
b[64619] == 64619 && 
b[64620] == 64620 && 
b[64621] == 64621 && 
b[64622] == 64622 && 
b[64623] == 64623 && 
b[64624] == 64624 && 
b[64625] == 64625 && 
b[64626] == 64626 && 
b[64627] == 64627 && 
b[64628] == 64628 && 
b[64629] == 64629 && 
b[64630] == 64630 && 
b[64631] == 64631 && 
b[64632] == 64632 && 
b[64633] == 64633 && 
b[64634] == 64634 && 
b[64635] == 64635 && 
b[64636] == 64636 && 
b[64637] == 64637 && 
b[64638] == 64638 && 
b[64639] == 64639 && 
b[64640] == 64640 && 
b[64641] == 64641 && 
b[64642] == 64642 && 
b[64643] == 64643 && 
b[64644] == 64644 && 
b[64645] == 64645 && 
b[64646] == 64646 && 
b[64647] == 64647 && 
b[64648] == 64648 && 
b[64649] == 64649 && 
b[64650] == 64650 && 
b[64651] == 64651 && 
b[64652] == 64652 && 
b[64653] == 64653 && 
b[64654] == 64654 && 
b[64655] == 64655 && 
b[64656] == 64656 && 
b[64657] == 64657 && 
b[64658] == 64658 && 
b[64659] == 64659 && 
b[64660] == 64660 && 
b[64661] == 64661 && 
b[64662] == 64662 && 
b[64663] == 64663 && 
b[64664] == 64664 && 
b[64665] == 64665 && 
b[64666] == 64666 && 
b[64667] == 64667 && 
b[64668] == 64668 && 
b[64669] == 64669 && 
b[64670] == 64670 && 
b[64671] == 64671 && 
b[64672] == 64672 && 
b[64673] == 64673 && 
b[64674] == 64674 && 
b[64675] == 64675 && 
b[64676] == 64676 && 
b[64677] == 64677 && 
b[64678] == 64678 && 
b[64679] == 64679 && 
b[64680] == 64680 && 
b[64681] == 64681 && 
b[64682] == 64682 && 
b[64683] == 64683 && 
b[64684] == 64684 && 
b[64685] == 64685 && 
b[64686] == 64686 && 
b[64687] == 64687 && 
b[64688] == 64688 && 
b[64689] == 64689 && 
b[64690] == 64690 && 
b[64691] == 64691 && 
b[64692] == 64692 && 
b[64693] == 64693 && 
b[64694] == 64694 && 
b[64695] == 64695 && 
b[64696] == 64696 && 
b[64697] == 64697 && 
b[64698] == 64698 && 
b[64699] == 64699 && 
b[64700] == 64700 && 
b[64701] == 64701 && 
b[64702] == 64702 && 
b[64703] == 64703 && 
b[64704] == 64704 && 
b[64705] == 64705 && 
b[64706] == 64706 && 
b[64707] == 64707 && 
b[64708] == 64708 && 
b[64709] == 64709 && 
b[64710] == 64710 && 
b[64711] == 64711 && 
b[64712] == 64712 && 
b[64713] == 64713 && 
b[64714] == 64714 && 
b[64715] == 64715 && 
b[64716] == 64716 && 
b[64717] == 64717 && 
b[64718] == 64718 && 
b[64719] == 64719 && 
b[64720] == 64720 && 
b[64721] == 64721 && 
b[64722] == 64722 && 
b[64723] == 64723 && 
b[64724] == 64724 && 
b[64725] == 64725 && 
b[64726] == 64726 && 
b[64727] == 64727 && 
b[64728] == 64728 && 
b[64729] == 64729 && 
b[64730] == 64730 && 
b[64731] == 64731 && 
b[64732] == 64732 && 
b[64733] == 64733 && 
b[64734] == 64734 && 
b[64735] == 64735 && 
b[64736] == 64736 && 
b[64737] == 64737 && 
b[64738] == 64738 && 
b[64739] == 64739 && 
b[64740] == 64740 && 
b[64741] == 64741 && 
b[64742] == 64742 && 
b[64743] == 64743 && 
b[64744] == 64744 && 
b[64745] == 64745 && 
b[64746] == 64746 && 
b[64747] == 64747 && 
b[64748] == 64748 && 
b[64749] == 64749 && 
b[64750] == 64750 && 
b[64751] == 64751 && 
b[64752] == 64752 && 
b[64753] == 64753 && 
b[64754] == 64754 && 
b[64755] == 64755 && 
b[64756] == 64756 && 
b[64757] == 64757 && 
b[64758] == 64758 && 
b[64759] == 64759 && 
b[64760] == 64760 && 
b[64761] == 64761 && 
b[64762] == 64762 && 
b[64763] == 64763 && 
b[64764] == 64764 && 
b[64765] == 64765 && 
b[64766] == 64766 && 
b[64767] == 64767 && 
b[64768] == 64768 && 
b[64769] == 64769 && 
b[64770] == 64770 && 
b[64771] == 64771 && 
b[64772] == 64772 && 
b[64773] == 64773 && 
b[64774] == 64774 && 
b[64775] == 64775 && 
b[64776] == 64776 && 
b[64777] == 64777 && 
b[64778] == 64778 && 
b[64779] == 64779 && 
b[64780] == 64780 && 
b[64781] == 64781 && 
b[64782] == 64782 && 
b[64783] == 64783 && 
b[64784] == 64784 && 
b[64785] == 64785 && 
b[64786] == 64786 && 
b[64787] == 64787 && 
b[64788] == 64788 && 
b[64789] == 64789 && 
b[64790] == 64790 && 
b[64791] == 64791 && 
b[64792] == 64792 && 
b[64793] == 64793 && 
b[64794] == 64794 && 
b[64795] == 64795 && 
b[64796] == 64796 && 
b[64797] == 64797 && 
b[64798] == 64798 && 
b[64799] == 64799 && 
b[64800] == 64800 && 
b[64801] == 64801 && 
b[64802] == 64802 && 
b[64803] == 64803 && 
b[64804] == 64804 && 
b[64805] == 64805 && 
b[64806] == 64806 && 
b[64807] == 64807 && 
b[64808] == 64808 && 
b[64809] == 64809 && 
b[64810] == 64810 && 
b[64811] == 64811 && 
b[64812] == 64812 && 
b[64813] == 64813 && 
b[64814] == 64814 && 
b[64815] == 64815 && 
b[64816] == 64816 && 
b[64817] == 64817 && 
b[64818] == 64818 && 
b[64819] == 64819 && 
b[64820] == 64820 && 
b[64821] == 64821 && 
b[64822] == 64822 && 
b[64823] == 64823 && 
b[64824] == 64824 && 
b[64825] == 64825 && 
b[64826] == 64826 && 
b[64827] == 64827 && 
b[64828] == 64828 && 
b[64829] == 64829 && 
b[64830] == 64830 && 
b[64831] == 64831 && 
b[64832] == 64832 && 
b[64833] == 64833 && 
b[64834] == 64834 && 
b[64835] == 64835 && 
b[64836] == 64836 && 
b[64837] == 64837 && 
b[64838] == 64838 && 
b[64839] == 64839 && 
b[64840] == 64840 && 
b[64841] == 64841 && 
b[64842] == 64842 && 
b[64843] == 64843 && 
b[64844] == 64844 && 
b[64845] == 64845 && 
b[64846] == 64846 && 
b[64847] == 64847 && 
b[64848] == 64848 && 
b[64849] == 64849 && 
b[64850] == 64850 && 
b[64851] == 64851 && 
b[64852] == 64852 && 
b[64853] == 64853 && 
b[64854] == 64854 && 
b[64855] == 64855 && 
b[64856] == 64856 && 
b[64857] == 64857 && 
b[64858] == 64858 && 
b[64859] == 64859 && 
b[64860] == 64860 && 
b[64861] == 64861 && 
b[64862] == 64862 && 
b[64863] == 64863 && 
b[64864] == 64864 && 
b[64865] == 64865 && 
b[64866] == 64866 && 
b[64867] == 64867 && 
b[64868] == 64868 && 
b[64869] == 64869 && 
b[64870] == 64870 && 
b[64871] == 64871 && 
b[64872] == 64872 && 
b[64873] == 64873 && 
b[64874] == 64874 && 
b[64875] == 64875 && 
b[64876] == 64876 && 
b[64877] == 64877 && 
b[64878] == 64878 && 
b[64879] == 64879 && 
b[64880] == 64880 && 
b[64881] == 64881 && 
b[64882] == 64882 && 
b[64883] == 64883 && 
b[64884] == 64884 && 
b[64885] == 64885 && 
b[64886] == 64886 && 
b[64887] == 64887 && 
b[64888] == 64888 && 
b[64889] == 64889 && 
b[64890] == 64890 && 
b[64891] == 64891 && 
b[64892] == 64892 && 
b[64893] == 64893 && 
b[64894] == 64894 && 
b[64895] == 64895 && 
b[64896] == 64896 && 
b[64897] == 64897 && 
b[64898] == 64898 && 
b[64899] == 64899 && 
b[64900] == 64900 && 
b[64901] == 64901 && 
b[64902] == 64902 && 
b[64903] == 64903 && 
b[64904] == 64904 && 
b[64905] == 64905 && 
b[64906] == 64906 && 
b[64907] == 64907 && 
b[64908] == 64908 && 
b[64909] == 64909 && 
b[64910] == 64910 && 
b[64911] == 64911 && 
b[64912] == 64912 && 
b[64913] == 64913 && 
b[64914] == 64914 && 
b[64915] == 64915 && 
b[64916] == 64916 && 
b[64917] == 64917 && 
b[64918] == 64918 && 
b[64919] == 64919 && 
b[64920] == 64920 && 
b[64921] == 64921 && 
b[64922] == 64922 && 
b[64923] == 64923 && 
b[64924] == 64924 && 
b[64925] == 64925 && 
b[64926] == 64926 && 
b[64927] == 64927 && 
b[64928] == 64928 && 
b[64929] == 64929 && 
b[64930] == 64930 && 
b[64931] == 64931 && 
b[64932] == 64932 && 
b[64933] == 64933 && 
b[64934] == 64934 && 
b[64935] == 64935 && 
b[64936] == 64936 && 
b[64937] == 64937 && 
b[64938] == 64938 && 
b[64939] == 64939 && 
b[64940] == 64940 && 
b[64941] == 64941 && 
b[64942] == 64942 && 
b[64943] == 64943 && 
b[64944] == 64944 && 
b[64945] == 64945 && 
b[64946] == 64946 && 
b[64947] == 64947 && 
b[64948] == 64948 && 
b[64949] == 64949 && 
b[64950] == 64950 && 
b[64951] == 64951 && 
b[64952] == 64952 && 
b[64953] == 64953 && 
b[64954] == 64954 && 
b[64955] == 64955 && 
b[64956] == 64956 && 
b[64957] == 64957 && 
b[64958] == 64958 && 
b[64959] == 64959 && 
b[64960] == 64960 && 
b[64961] == 64961 && 
b[64962] == 64962 && 
b[64963] == 64963 && 
b[64964] == 64964 && 
b[64965] == 64965 && 
b[64966] == 64966 && 
b[64967] == 64967 && 
b[64968] == 64968 && 
b[64969] == 64969 && 
b[64970] == 64970 && 
b[64971] == 64971 && 
b[64972] == 64972 && 
b[64973] == 64973 && 
b[64974] == 64974 && 
b[64975] == 64975 && 
b[64976] == 64976 && 
b[64977] == 64977 && 
b[64978] == 64978 && 
b[64979] == 64979 && 
b[64980] == 64980 && 
b[64981] == 64981 && 
b[64982] == 64982 && 
b[64983] == 64983 && 
b[64984] == 64984 && 
b[64985] == 64985 && 
b[64986] == 64986 && 
b[64987] == 64987 && 
b[64988] == 64988 && 
b[64989] == 64989 && 
b[64990] == 64990 && 
b[64991] == 64991 && 
b[64992] == 64992 && 
b[64993] == 64993 && 
b[64994] == 64994 && 
b[64995] == 64995 && 
b[64996] == 64996 && 
b[64997] == 64997 && 
b[64998] == 64998 && 
b[64999] == 64999 && 
b[65000] == 65000 && 
b[65001] == 65001 && 
b[65002] == 65002 && 
b[65003] == 65003 && 
b[65004] == 65004 && 
b[65005] == 65005 && 
b[65006] == 65006 && 
b[65007] == 65007 && 
b[65008] == 65008 && 
b[65009] == 65009 && 
b[65010] == 65010 && 
b[65011] == 65011 && 
b[65012] == 65012 && 
b[65013] == 65013 && 
b[65014] == 65014 && 
b[65015] == 65015 && 
b[65016] == 65016 && 
b[65017] == 65017 && 
b[65018] == 65018 && 
b[65019] == 65019 && 
b[65020] == 65020 && 
b[65021] == 65021 && 
b[65022] == 65022 && 
b[65023] == 65023 && 
b[65024] == 65024 && 
b[65025] == 65025 && 
b[65026] == 65026 && 
b[65027] == 65027 && 
b[65028] == 65028 && 
b[65029] == 65029 && 
b[65030] == 65030 && 
b[65031] == 65031 && 
b[65032] == 65032 && 
b[65033] == 65033 && 
b[65034] == 65034 && 
b[65035] == 65035 && 
b[65036] == 65036 && 
b[65037] == 65037 && 
b[65038] == 65038 && 
b[65039] == 65039 && 
b[65040] == 65040 && 
b[65041] == 65041 && 
b[65042] == 65042 && 
b[65043] == 65043 && 
b[65044] == 65044 && 
b[65045] == 65045 && 
b[65046] == 65046 && 
b[65047] == 65047 && 
b[65048] == 65048 && 
b[65049] == 65049 && 
b[65050] == 65050 && 
b[65051] == 65051 && 
b[65052] == 65052 && 
b[65053] == 65053 && 
b[65054] == 65054 && 
b[65055] == 65055 && 
b[65056] == 65056 && 
b[65057] == 65057 && 
b[65058] == 65058 && 
b[65059] == 65059 && 
b[65060] == 65060 && 
b[65061] == 65061 && 
b[65062] == 65062 && 
b[65063] == 65063 && 
b[65064] == 65064 && 
b[65065] == 65065 && 
b[65066] == 65066 && 
b[65067] == 65067 && 
b[65068] == 65068 && 
b[65069] == 65069 && 
b[65070] == 65070 && 
b[65071] == 65071 && 
b[65072] == 65072 && 
b[65073] == 65073 && 
b[65074] == 65074 && 
b[65075] == 65075 && 
b[65076] == 65076 && 
b[65077] == 65077 && 
b[65078] == 65078 && 
b[65079] == 65079 && 
b[65080] == 65080 && 
b[65081] == 65081 && 
b[65082] == 65082 && 
b[65083] == 65083 && 
b[65084] == 65084 && 
b[65085] == 65085 && 
b[65086] == 65086 && 
b[65087] == 65087 && 
b[65088] == 65088 && 
b[65089] == 65089 && 
b[65090] == 65090 && 
b[65091] == 65091 && 
b[65092] == 65092 && 
b[65093] == 65093 && 
b[65094] == 65094 && 
b[65095] == 65095 && 
b[65096] == 65096 && 
b[65097] == 65097 && 
b[65098] == 65098 && 
b[65099] == 65099 && 
b[65100] == 65100 && 
b[65101] == 65101 && 
b[65102] == 65102 && 
b[65103] == 65103 && 
b[65104] == 65104 && 
b[65105] == 65105 && 
b[65106] == 65106 && 
b[65107] == 65107 && 
b[65108] == 65108 && 
b[65109] == 65109 && 
b[65110] == 65110 && 
b[65111] == 65111 && 
b[65112] == 65112 && 
b[65113] == 65113 && 
b[65114] == 65114 && 
b[65115] == 65115 && 
b[65116] == 65116 && 
b[65117] == 65117 && 
b[65118] == 65118 && 
b[65119] == 65119 && 
b[65120] == 65120 && 
b[65121] == 65121 && 
b[65122] == 65122 && 
b[65123] == 65123 && 
b[65124] == 65124 && 
b[65125] == 65125 && 
b[65126] == 65126 && 
b[65127] == 65127 && 
b[65128] == 65128 && 
b[65129] == 65129 && 
b[65130] == 65130 && 
b[65131] == 65131 && 
b[65132] == 65132 && 
b[65133] == 65133 && 
b[65134] == 65134 && 
b[65135] == 65135 && 
b[65136] == 65136 && 
b[65137] == 65137 && 
b[65138] == 65138 && 
b[65139] == 65139 && 
b[65140] == 65140 && 
b[65141] == 65141 && 
b[65142] == 65142 && 
b[65143] == 65143 && 
b[65144] == 65144 && 
b[65145] == 65145 && 
b[65146] == 65146 && 
b[65147] == 65147 && 
b[65148] == 65148 && 
b[65149] == 65149 && 
b[65150] == 65150 && 
b[65151] == 65151 && 
b[65152] == 65152 && 
b[65153] == 65153 && 
b[65154] == 65154 && 
b[65155] == 65155 && 
b[65156] == 65156 && 
b[65157] == 65157 && 
b[65158] == 65158 && 
b[65159] == 65159 && 
b[65160] == 65160 && 
b[65161] == 65161 && 
b[65162] == 65162 && 
b[65163] == 65163 && 
b[65164] == 65164 && 
b[65165] == 65165 && 
b[65166] == 65166 && 
b[65167] == 65167 && 
b[65168] == 65168 && 
b[65169] == 65169 && 
b[65170] == 65170 && 
b[65171] == 65171 && 
b[65172] == 65172 && 
b[65173] == 65173 && 
b[65174] == 65174 && 
b[65175] == 65175 && 
b[65176] == 65176 && 
b[65177] == 65177 && 
b[65178] == 65178 && 
b[65179] == 65179 && 
b[65180] == 65180 && 
b[65181] == 65181 && 
b[65182] == 65182 && 
b[65183] == 65183 && 
b[65184] == 65184 && 
b[65185] == 65185 && 
b[65186] == 65186 && 
b[65187] == 65187 && 
b[65188] == 65188 && 
b[65189] == 65189 && 
b[65190] == 65190 && 
b[65191] == 65191 && 
b[65192] == 65192 && 
b[65193] == 65193 && 
b[65194] == 65194 && 
b[65195] == 65195 && 
b[65196] == 65196 && 
b[65197] == 65197 && 
b[65198] == 65198 && 
b[65199] == 65199 && 
b[65200] == 65200 && 
b[65201] == 65201 && 
b[65202] == 65202 && 
b[65203] == 65203 && 
b[65204] == 65204 && 
b[65205] == 65205 && 
b[65206] == 65206 && 
b[65207] == 65207 && 
b[65208] == 65208 && 
b[65209] == 65209 && 
b[65210] == 65210 && 
b[65211] == 65211 && 
b[65212] == 65212 && 
b[65213] == 65213 && 
b[65214] == 65214 && 
b[65215] == 65215 && 
b[65216] == 65216 && 
b[65217] == 65217 && 
b[65218] == 65218 && 
b[65219] == 65219 && 
b[65220] == 65220 && 
b[65221] == 65221 && 
b[65222] == 65222 && 
b[65223] == 65223 && 
b[65224] == 65224 && 
b[65225] == 65225 && 
b[65226] == 65226 && 
b[65227] == 65227 && 
b[65228] == 65228 && 
b[65229] == 65229 && 
b[65230] == 65230 && 
b[65231] == 65231 && 
b[65232] == 65232 && 
b[65233] == 65233 && 
b[65234] == 65234 && 
b[65235] == 65235 && 
b[65236] == 65236 && 
b[65237] == 65237 && 
b[65238] == 65238 && 
b[65239] == 65239 && 
b[65240] == 65240 && 
b[65241] == 65241 && 
b[65242] == 65242 && 
b[65243] == 65243 && 
b[65244] == 65244 && 
b[65245] == 65245 && 
b[65246] == 65246 && 
b[65247] == 65247 && 
b[65248] == 65248 && 
b[65249] == 65249 && 
b[65250] == 65250 && 
b[65251] == 65251 && 
b[65252] == 65252 && 
b[65253] == 65253 && 
b[65254] == 65254 && 
b[65255] == 65255 && 
b[65256] == 65256 && 
b[65257] == 65257 && 
b[65258] == 65258 && 
b[65259] == 65259 && 
b[65260] == 65260 && 
b[65261] == 65261 && 
b[65262] == 65262 && 
b[65263] == 65263 && 
b[65264] == 65264 && 
b[65265] == 65265 && 
b[65266] == 65266 && 
b[65267] == 65267 && 
b[65268] == 65268 && 
b[65269] == 65269 && 
b[65270] == 65270 && 
b[65271] == 65271 && 
b[65272] == 65272 && 
b[65273] == 65273 && 
b[65274] == 65274 && 
b[65275] == 65275 && 
b[65276] == 65276 && 
b[65277] == 65277 && 
b[65278] == 65278 && 
b[65279] == 65279 && 
b[65280] == 65280 && 
b[65281] == 65281 && 
b[65282] == 65282 && 
b[65283] == 65283 && 
b[65284] == 65284 && 
b[65285] == 65285 && 
b[65286] == 65286 && 
b[65287] == 65287 && 
b[65288] == 65288 && 
b[65289] == 65289 && 
b[65290] == 65290 && 
b[65291] == 65291 && 
b[65292] == 65292 && 
b[65293] == 65293 && 
b[65294] == 65294 && 
b[65295] == 65295 && 
b[65296] == 65296 && 
b[65297] == 65297 && 
b[65298] == 65298 && 
b[65299] == 65299 && 
b[65300] == 65300 && 
b[65301] == 65301 && 
b[65302] == 65302 && 
b[65303] == 65303 && 
b[65304] == 65304 && 
b[65305] == 65305 && 
b[65306] == 65306 && 
b[65307] == 65307 && 
b[65308] == 65308 && 
b[65309] == 65309 && 
b[65310] == 65310 && 
b[65311] == 65311 && 
b[65312] == 65312 && 
b[65313] == 65313 && 
b[65314] == 65314 && 
b[65315] == 65315 && 
b[65316] == 65316 && 
b[65317] == 65317 && 
b[65318] == 65318 && 
b[65319] == 65319 && 
b[65320] == 65320 && 
b[65321] == 65321 && 
b[65322] == 65322 && 
b[65323] == 65323 && 
b[65324] == 65324 && 
b[65325] == 65325 && 
b[65326] == 65326 && 
b[65327] == 65327 && 
b[65328] == 65328 && 
b[65329] == 65329 && 
b[65330] == 65330 && 
b[65331] == 65331 && 
b[65332] == 65332 && 
b[65333] == 65333 && 
b[65334] == 65334 && 
b[65335] == 65335 && 
b[65336] == 65336 && 
b[65337] == 65337 && 
b[65338] == 65338 && 
b[65339] == 65339 && 
b[65340] == 65340 && 
b[65341] == 65341 && 
b[65342] == 65342 && 
b[65343] == 65343 && 
b[65344] == 65344 && 
b[65345] == 65345 && 
b[65346] == 65346 && 
b[65347] == 65347 && 
b[65348] == 65348 && 
b[65349] == 65349 && 
b[65350] == 65350 && 
b[65351] == 65351 && 
b[65352] == 65352 && 
b[65353] == 65353 && 
b[65354] == 65354 && 
b[65355] == 65355 && 
b[65356] == 65356 && 
b[65357] == 65357 && 
b[65358] == 65358 && 
b[65359] == 65359 && 
b[65360] == 65360 && 
b[65361] == 65361 && 
b[65362] == 65362 && 
b[65363] == 65363 && 
b[65364] == 65364 && 
b[65365] == 65365 && 
b[65366] == 65366 && 
b[65367] == 65367 && 
b[65368] == 65368 && 
b[65369] == 65369 && 
b[65370] == 65370 && 
b[65371] == 65371 && 
b[65372] == 65372 && 
b[65373] == 65373 && 
b[65374] == 65374 && 
b[65375] == 65375 && 
b[65376] == 65376 && 
b[65377] == 65377 && 
b[65378] == 65378 && 
b[65379] == 65379 && 
b[65380] == 65380 && 
b[65381] == 65381 && 
b[65382] == 65382 && 
b[65383] == 65383 && 
b[65384] == 65384 && 
b[65385] == 65385 && 
b[65386] == 65386 && 
b[65387] == 65387 && 
b[65388] == 65388 && 
b[65389] == 65389 && 
b[65390] == 65390 && 
b[65391] == 65391 && 
b[65392] == 65392 && 
b[65393] == 65393 && 
b[65394] == 65394 && 
b[65395] == 65395 && 
b[65396] == 65396 && 
b[65397] == 65397 && 
b[65398] == 65398 && 
b[65399] == 65399 && 
b[65400] == 65400 && 
b[65401] == 65401 && 
b[65402] == 65402 && 
b[65403] == 65403 && 
b[65404] == 65404 && 
b[65405] == 65405 && 
b[65406] == 65406 && 
b[65407] == 65407 && 
b[65408] == 65408 && 
b[65409] == 65409 && 
b[65410] == 65410 && 
b[65411] == 65411 && 
b[65412] == 65412 && 
b[65413] == 65413 && 
b[65414] == 65414 && 
b[65415] == 65415 && 
b[65416] == 65416 && 
b[65417] == 65417 && 
b[65418] == 65418 && 
b[65419] == 65419 && 
b[65420] == 65420 && 
b[65421] == 65421 && 
b[65422] == 65422 && 
b[65423] == 65423 && 
b[65424] == 65424 && 
b[65425] == 65425 && 
b[65426] == 65426 && 
b[65427] == 65427 && 
b[65428] == 65428 && 
b[65429] == 65429 && 
b[65430] == 65430 && 
b[65431] == 65431 && 
b[65432] == 65432 && 
b[65433] == 65433 && 
b[65434] == 65434 && 
b[65435] == 65435 && 
b[65436] == 65436 && 
b[65437] == 65437 && 
b[65438] == 65438 && 
b[65439] == 65439 && 
b[65440] == 65440 && 
b[65441] == 65441 && 
b[65442] == 65442 && 
b[65443] == 65443 && 
b[65444] == 65444 && 
b[65445] == 65445 && 
b[65446] == 65446 && 
b[65447] == 65447 && 
b[65448] == 65448 && 
b[65449] == 65449 && 
b[65450] == 65450 && 
b[65451] == 65451 && 
b[65452] == 65452 && 
b[65453] == 65453 && 
b[65454] == 65454 && 
b[65455] == 65455 && 
b[65456] == 65456 && 
b[65457] == 65457 && 
b[65458] == 65458 && 
b[65459] == 65459 && 
b[65460] == 65460 && 
b[65461] == 65461 && 
b[65462] == 65462 && 
b[65463] == 65463 && 
b[65464] == 65464 && 
b[65465] == 65465 && 
b[65466] == 65466 && 
b[65467] == 65467 && 
b[65468] == 65468 && 
b[65469] == 65469 && 
b[65470] == 65470 && 
b[65471] == 65471 && 
b[65472] == 65472 && 
b[65473] == 65473 && 
b[65474] == 65474 && 
b[65475] == 65475 && 
b[65476] == 65476 && 
b[65477] == 65477 && 
b[65478] == 65478 && 
b[65479] == 65479 && 
b[65480] == 65480 && 
b[65481] == 65481 && 
b[65482] == 65482 && 
b[65483] == 65483 && 
b[65484] == 65484 && 
b[65485] == 65485 && 
b[65486] == 65486 && 
b[65487] == 65487 && 
b[65488] == 65488 && 
b[65489] == 65489 && 
b[65490] == 65490 && 
b[65491] == 65491 && 
b[65492] == 65492 && 
b[65493] == 65493 && 
b[65494] == 65494 && 
b[65495] == 65495 && 
b[65496] == 65496 && 
b[65497] == 65497 && 
b[65498] == 65498 && 
b[65499] == 65499 && 
b[65500] == 65500 && 
b[65501] == 65501 && 
b[65502] == 65502 && 
b[65503] == 65503 && 
b[65504] == 65504 && 
b[65505] == 65505 && 
b[65506] == 65506 && 
b[65507] == 65507 && 
b[65508] == 65508 && 
b[65509] == 65509 && 
b[65510] == 65510 && 
b[65511] == 65511 && 
b[65512] == 65512 && 
b[65513] == 65513 && 
b[65514] == 65514 && 
b[65515] == 65515 && 
b[65516] == 65516 && 
b[65517] == 65517 && 
b[65518] == 65518 && 
b[65519] == 65519 && 
b[65520] == 65520 && 
b[65521] == 65521 && 
b[65522] == 65522 && 
b[65523] == 65523 && 
b[65524] == 65524 && 
b[65525] == 65525 && 
b[65526] == 65526 && 
b[65527] == 65527 && 
b[65528] == 65528 && 
b[65529] == 65529 && 
b[65530] == 65530 && 
b[65531] == 65531 && 
b[65532] == 65532 && 
b[65533] == 65533 && 
b[65534] == 65534 && 
b[65535] == 65535 
));

//G(parity=0);

endmodule // slidingBoard
